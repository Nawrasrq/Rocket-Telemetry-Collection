PK   ���X_d�y  H�     cirkitFile.json�]m�۸��+S�/wU�B��|�nrWn��l���k
$�]diBQ~���=J�%����h.wS����n4���~�T�[����t�z�ZNn��NLe?�ç�t�8_�׫��*��0�����/�.*VWK���cWh�5�d��N�(���D�i%���.��'���O�����9�] {3Ks+��GqV��lY��(X�*+��2��wVl�˔t<F�H�LG��6JYɔ�.��O�yy�3^�8�*w�d"��yTz.e��Y
JZ,i�(��:�w�&\��Ņ�zKg��I���Rk-�K�L譄�ٺ��Q�3��)M�h�6�hT��xR�n��f�"���TF��=��]�ǌ��L9#�B���D��4��8�q�s�4�T߁�<pA�'��ǉ��D�q"�8"�[_�5��#��E2���Ħ�t�HX[K���
JՌRu��C1�5��E�%�EL*���Q���\Y&S�Ta{����5c{�Pu߂��	�꾅��}�F�'�FSj&�����o�Q����oБ���X�ABzp�����r �� ��Hc���0(�~���� d�Us��L\�� ��KLQl�t�9:Q���ӌ��@���'δ�P�O�0�����F�&.1m�)�K�d��f
�"��eG�K/�fdP���������P3���>P�Z�*�>�����;���
 ��"��\�� �� R� R��R�1#II�蒅A] ��A/��W�\R�4��K�Ҵ	`�,��#&�Y�0(�lp#�E1aP�à��A1�b�<�E�l	6fD���f��m6�@>�1�|��(as�þ6O@�QC�M��2jf���a�`s��x��g�[����2:�؜m )�#�������FlR6�.��	6�:<�)� S`ܯG'AC�	��q��!f�#B�IC�	�q��<��<��T��4�h4��M5�Mg3�)�a?��۷�95��M����ԕYSst)<�D�"E�����HI�H� .xà���/�_�,�Y�0fa@� ��A1d�à��A1�b�<�y�0(�aP, X�����K	���B����Sst)���N�ѥ��Q3�N�ѥ�tj�.et�ѩ9��ёF���RFG���K]MЩ9��ѵ�� &z��z|j.��0 ��� b�`xܯǧ�ŠSst)�F���RF�N�ѥ��mlj�.�P�oS���z{f�~n?OnY:�|�Wn}��0����������ܾ��У$��O)�����kUݼ�Ey���\�մ�I��u8�`%�f��R}5S^�ǟG'g'yl=uS�E��@z���Q����_�fd�@i
�i��72mr���o ���fB�ܔ��5�z�R3�ަ��\b�@���r�/Ĺ�kr��ֺHc�h�L#���ʠ�Q�mU��R�mFqS�P�W3rn����r��2�{{�z?��D��3����A���㌽d��S6�rV��7KەYy:q��WK�4
|?\z�g�+�Az���!v�	��#]�|Z��5E���뱞F�t���r��� ���uM�Q�E�v��L�nP����b*��1�w1��=:
��=zC6�DL>��I/�n�.�������yl^"�J� 1�z�!x�Y@���R �G��Z�M
_�)��/�`Sį{5x�T��`��X*����a�g�.���rp�uI�@�{��/���uIΝ�� �Kfj�CA]�
��� �0X �8]lY�n<],k����l@oC�
�0< ��Jz?���n���E��We����R��[����"��������CI�K�:�Tڮ&M}�N�uD_P@Q'����V*\���z�g��o$8�G�|�
���%� *f��H�0eT�r*N9٬R�js� I ���DNE"�"�S�ȩHl�8�/č�y���Q��֮��S�ft���ϫ�/8G٥��;Jbc� �/����G�AقN��<�
��֡/���.��
���/��wg��C�3@Q'E�]�U8����!/� I �C~:������ I��w��L�G ����	�`��X 7��7�L���v�;���d*З���X6��#q����Y���d�_�lƗ���Ω�(�@���p�����{���k>��<e�����3O�<5����3��<����9�����{�9�����9����~��͞����?�
��`��%;T�L���`���7���f���=���;'��X�+Nc&���i��O�!}��v
��P,5���IJ��(A�	%��:��W�)�)ŵ'��:���I�J�F:-p�	}�}���e4�{����e������ke�o�Z��-��d�����7~N�����]�8-��"yZ�vE괈��iQ�+JN���H�����Q5��}^9c������~1_�[d���?���|_�Go�գ���ޮ�1�����-f"���)K�,�R���IA��7��L��D,d�4��4�R�Uz�%�q췹���uS�N�ͮͲ�
By��ɪ���Us�y���U�p���K���)�����MQ�p��g�$V��j7ܻr��`(��Y����A\:K25�<����X��.?(�y�K���վ�6�������ɇǥ���$P��j��Z�4��t:�h���&x�l�s�	�k������G�;�-�b�p�_��y�p�g���f^9���8�f�)MQo*W)pHv����B Mڀ�Х���V��"��+�H+p�q �y���h���(���:ҸNf�P�d�U����a�D��&8N��IS8i	NZ��&���T��d�_��� _���9o��i�_���G{:�qt���M�h]�����	��'8R���zʔ�/k�S�%�e[����>9���� �)�:�U�z�����u���]c��&�w���\]<�M�w��m��^gDĔ4��Z�D���'e�Db]bz��q�3�����͖�ۜ�T%��-,��i�s�RZ��<˜ix}�|�KS�?���k�T��,�X3�Y	�t��f�����,82JҸ��GE�����F�D�E�m����΋�	���iynɏ�=���̬6)88�FE&�!3��>.�VW�h�jU���RR��.A?���6s�Fe���Ɖ��vH�q�Z�Cm�ɕ��F�qmX�O�(��e�Le������h��y>�(³������ϗ[�ۇ��cu�Y��C¿<����om���]ٷ)�J�i9_�p��;�O �TE0� ��q�0^���)˓2�} +�ԘȔ�/䥆X|:U� �g�`%�u������dY�ť��)mfEb���L�,s�"k\���#?�Q�gE��T����z7���ۛ��7���7_��77���Tw�e���%7����UnzS�n���fN�-P�߶5��U��f��S�Ggjg_�m5��-\Q7�i��6������/�m;U���tao�A(�\Uk�j3�o�,���@KB��2�h�����x�T�Nl�X"��\s���De��H�E�\�f�j܉E�菝X���<qc%�"j*��e�?>ޑ��:X��j|%�n${z~�O��Q��	}Ġ�
~ܱ�-�����*��2ɲ�^ft-E+�/�L�(#�9��Hf!��e��4�ىG.jc�\%=r��/6��z���s�m�N�Z�{�n�!�o=O�-�j���s���l���LҝR��Nu�:iQ'�ItRɮ�ߔ�0�)c�ED
3V��D�i,���t� Vj�(Q=t��$U��S`R�,���5����O���3���-�N:�$�!vmH�����$�J�|�S*0^)i���c���  �g���%U3�c!�kIkB관@D���H�<�Ҕ9��N���Ț��	��&��Cv`j�$�NR�0�d�9�#c1gC:c c���]��d���!�%L�L�+0�v_�5Xp{�L ��n"	1���a6bgp�.E��R�O�ϐI �.���<Y���bv��:r����>�U|&Y�U�{"_ >*}�y	�!�ۥ%Kvs{*�.۾�T-%Υ��:�¼� &t�����L��9�C�8Z��>�#�R��ެo���~�G��qYm��AJ���Dj������O��؜��4�����d6������{�I��?�~i����L����=�����/��ݧ��w���>����	hw��n�H�Ԫ~;_����?&����vP�J#�2�~	��c8�W�e����,���&~����/����k���������o�~�_=���J"qO���c$U{�kO���C�������@��σ( @qP ��Pk��@GT���i������n����@ۺH���;�?
�3�;>�ݽ��&�~0����N0ک $�<�R���s���]���w��Z�8C�+� ��S=�^�R�;�{-`�����1+I�H��s���"n!Af����0	^�3aqp ���󙸸?*�Q�#�g�S�zN�^*va8d�N�6�3ԣ�=�*�v+�VT����@�E,�_�̐/O\g���/��\z�k�E������E`��ic�P���9c��ٳ,4�xPs�H����M%ٱ{��-��X����uW���]�(��Q�vh���4�P��h�q�B�
	�\6�!�������}_ކ��6m*�:��9(�I�ځ�{��Z�8C�+�}I�ځ�{��Z�8C�+C��$����c�ݹ�n�n�������.#|Ƃs�j�2�ߵ�4�_?&;I�oc���
�j��Ȯe�O�z����n)tE�A���)ʮQ���T�a	���H�3,�)��b�s���]57����#e��2���?���,~X}xS��M�w�=��������[��qw�p��PK   ���Xx�آ  �  /   images/0fa89018-bbd7-413a-af56-bcf37033748d.png�b�PNG

   IHDR   d   V   9P3�   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  *IDATx��wl]Փ���ı��;�$!�З]B�e�!!�Z����X[ �(��Xjh�z
B'���q���W�|�y��ׅ��1�1ҳ���sϙ�9sf�;v�"r��Q4����OB��d2�A�pX��������Beee2h� �SPm�w����AZc1�F���lw���gͯ���'���J�$��СC���(�
����V����ѣGk�A5~O���M���� (�LJM]�̛T!w���ژD�!�%c��@�Yc' D�� &���J̡�f�$�J� 9�dڴi���k�HH�%�ɖ�[�8��cm2gB�������&�ׅ_Jk"������"��ƍS��ر#�x@����,---����Q�F����s��(�����e��s�g�J���=%�+��t�F#2n�U������TW׼��9眣���#�t������Ν;{Q�,���q����G���D'���J<��3��#O��\j��U��D2%sgM�yN�x�6�.�U{�HA}}�^�1j
p`=z����D��;}oj���


��2~C:<�@<�:oy<nj�r�D�FP'���xO)�J��c����Y�ُ���&�]�k���R9�/GHqa�4��p�;���TR��OQ��E\���㠃�M�6�y��db��0����WF���K
0t�gȤI�䭷ޒ�7�9� ^�l��^�Z+�s0,X X�����k�Icc�^�a��)S�s ��ɓe׮]
8����u��R��dZ��=E�>x������a\�;��΄�̊�
�6u�v�����}Q����v�y��d��@�nDR�N���uee�2��?Vi��_}��Jٺu�Ԍf����/�k��ʅ� �3�pHݬY��.����z�lu�m��#�Pp~��'-Ù�Z�/���V\II�����$۷oW��~����'� ��:�$262��$[��#�.�<�={�����|��r�7t� ��Y)����ŲaÆ�
���R�IW��t�I�xE/��dƌZ��ŋ�ꫯ�-[��ȑ#�1��\s�5RWW��P������'���=��	8�Ct,0$g���*Uo���p�M7i����ɦcЙ�������>�ߍ���rX�H�����t\J�c�jk��Eb)�u�2z�8�YWf.������혅
�1��=���Çk/E�ظ�� 'NTFқ� ���3g�|��Za: ���)�zP*ꩧ�R�2�Db�>$�:�l����7o��"�^�����UR�����${�w�R[�*��������:�*<q��)�g���u;!��
�� ��3OQ/=���F��7�Ș1c��W_�?�P�����2w�\�Ρ?C>�`w  ����`���OhYH��T!MH�������߫� ��~���By��������˵��N�!�0�Fh������Q��'�DNB���)�؛9`��i�����ʤ�$�7���8Go��w�;ϢWb��a���8Gg���Yc<�c�1Á�%v���y���`?�f��A�w�|�f BŹ���7d�Y�@���{~y���ٝO~�y��=6����<�v�>�����5��@��h��V@  	��_Ȍ�}A�f*��eo��s�.�R�jh���3H���3�����[�N�*}��eȐ!q�4;F���a�t ���V�\�7����}���g��=;���k�������:��h�B�vn�����+������[Z�=R__�.-�N*��V7� ��_��{���l����F$�V+�9{��1&ӆ%��NbZ��y�%��__y�7�<`�� ���%�tx��kd����l�j
���I��y���-Z$�����X��D�K;�Ԙ#,]�TMG?n���@WY�.Ԯ�T�I���D�MGr��v7��<��꒒7�ٙ�PnA
p��1����u�D
��!��A�U_A����R�n�]��1
~���β�����N�@�F��p] �@WYQ�����đ��`��t}KB�w�J�mj�ۼ1[�B� �HI�jEX����z($�_���Z�}�a��ݚ�N!��ȧN��0s��1�L-��"�8�c���F�g�H�z �b<�p�MB��T;�t]�S�O�&�h�/��!�U�x�͍2���nc�t�j�J G'>�^�p�_�h�E�Ĺ3����Pi����(H���� ��d�S[AҰa�tn���q`����7��$!X�
'����g��'(�8%�*D��2p1+ʎ�h7A7�����J� ���O���O�s�N���z?�p'O�&9 R�jjk%�L8@
<E�^���$��MH���<����('��]x�r�w����JDM�t2�-X%' ĩDʣr�<����C���̘��vQ��Ia�С2u�Җ��o�%Mn��he8˪f{��@v�q>�cQ��I����!�|��w���W�X�Ki���.;d��p�PT}�P�E�wV��hHvn����~��<@��K.�D���kM�Aך�M�4��[^���[/���7��u�� ��]�s�YH�2��866�&L`�-�~ވ��:XY�l�dvr�s�@�$/��� �L<��e޼y��s��k)@�t�JD�ɪU�T@�}��&Lp=9_d���ى?��C�p0�$�ś�ER��x����#���tR�Ȕ��$�F���_�e>q` =F�YZ���<�TS*(K�,Q��>�leL!���3���` �H"��aB�O?�t�T R�,^��'�����娣��[n�Eˆ1䈑f�`�j!��I�ç�=�#%�c�~��3I��)^d�& �St'Y �"�o��0��=��)���=�\+GC��d<,lx�Vo��F���p�u��Ҋ�l�>��-S{��,�@���=CR�)0lĈ
,���V�0Yɠ!��z�6!�Z�%�����i$��y��B	E���"Ub�$�~��",�i�q\w饗�5�>I���䈑� ����$�����2��"�{  ��%#��9 �^$pPa��zc|��E}��Hׇ� �6n�$U;wHA8�ͺ�C�a0fӀ�{L�ӋmP �#1X3�ڀ�`^�/pY̜9SA`|���A�x.y^�w��u�Yr��kO��$/��b��{r���"��ޛ��Tz������ԛh�������E*S�2�"�Xs�3��'[^`A1�[Ќ���<]3ۿ��\/4����몺8O�Rb�����{UK 	 �9��*�sy�<#0zR�0�,4����ď�q\3a�SS)7!\�a��V"����eb�QYݨ�C���H����-���7"�0��PU��ެKT��٨],D �Ct;�H	����]W�}����M;�%��,���w��x�$Ԥͳ�UY�
p�H�!�[��Te�G!r��K&M�[��1z%!h�X<%�u���U7˟�gd���I���L�Bɔ<��/r����������ĤPJ���x �D C K��/~�Ie��as�\��W2��݊�Т�X<-����'����	�L�������+�5� �e�[�~�i�Rb��4az�Ԩa4��%ݭ�#D���L�2�j�?���GL.�3h�\:�*7��Q�*O~�NVn��1�C�Y��Glk���sp���������"�gT�ۛI%�i��2��^�"���rihIt��u���
�	���K�p�l7�_Is
��< H@B�	�J��ZJ���a��R��ܴ�(����c���=A��庽ݚ��x�9�sލ
�vi�5�텲���e�#%���'���0�`�m��{� p-�;ʲ}Q8G�|A1<��%����En�G�m��M���Z���~+����*q<)T�E:�x��u�����&HÒd�`=�5w �R }��u�2�� �o�@��܉'��Q��>�(�,�qm�> z��գj���ϒ	Σj���[��Z������ќ��GW~�˭��¹��L��A�2~�89z�Q���)���U�P(� ���\znWAz9q��֐���������ō� ��}��-NnLc&�}��w"t�G��K��id��1u���J��z▧cQ�	Rτ�P"��&���m��M�A��fI4g]��4y�	�:c�\����D+���Sϧ-[&�@����o@R� ���bׄLa �T��QI�x΄	t��T��~K`$�i ,�v� �����7߬ϥ ��$�D'�#P6φ���'�LK�̡2�x�;
���Qai���&����e�kO�NH��X(�z�� ������0�Wr���M��q?L<��<����%u�DٲG����!e0U��[il�� D։�j� �A"��`��ak�Xs���C��:H����,�8���F��7^��~�@��ր)����S����VC�@���[IH�t,�ض�@��'0����q �L��H	�[m �<��Q��'�z�\�h�m�a1v�D�%����8LjQ�n@{eo���霅I=������0ö����%�E"x�1a���r�e.gۆ�� �9�������~-�5�Ȳ� �&��vl�.���ݮ��裏�s�����W�Q��5`���{�����*b�~���1�����U=�2I�*�/7VuU6[�;��wk��R��������/>\"Sg�|�>vr`pF� -|�=���׸ep���v�m��Ʋ|� z�G�3_@uuLHd&|&��;ԭ�Z+������Z��0T��&��C9	aK���@�����xUF]�A�F`)inK���$�e�W�t�>s�`��'��A�i��E)�!m	�on�+[k(+�,�����̲�q��iji�������VI���-�Av����xf�����	e�dP��($� %DCa�<�Lj��6��D ���L�QW�.(&�~�r1�fϑ��BI�v��?�\%/}�IZڒ�#$�[��ѕ�x6���/|��Z�~�1����	��:3	�mn�D�ͻo'@pC�+΅�'��qeY?V8��b ��_�k�,[]3�7���kss�C~#4��X�~�㨓���oм洙������QS$R迫�� L��$�	��ф10.��F=Y�5a̳�>{5��Fi�Z��S�5�"�).w]p/^���pvi�@�9�3���x��'3t~[�pa�v��|�����w�G���_;�[kiy������Q��͒=�X������J���H��uQ"�񑁵go  `�$�n� ��ez���Q�|��ڵ�X_���?����i�rfN�[�!\�^t�Er뭷��%K�] �r�H&�ʮU���]""���j,�"���DVo�r�-����8�1��^#}�Q�%��8��$�X#���HVV0�B�f��z�v����%8KC�#�m\o	3�I5��Ww˨;d��Z�xp�n��[k0��6�[b������N�l��i�{��UW]��I"v`���n[k[f���{l�l�+ȼ�6�z���.���R��w��֨{CΖ� �J��!٬E�M �8�d��K�gk�MfI�0g0�;I�az^��?^N��1��%'�]��T r�P��00H�`5.D�-�X�3�r�0v�����"�$rP&�����I=�Y�ڣ�䘵����`N��e-8L$]���e[kpL��Z4�2a.�d�W&�0�,��~+�]B���=�\U+��}ѢEz��|�J�'xS9��=�7+,y@��z�ˍ����>��蝌aD-	�K �t�Ac|�X&]�!0]��G$�����L �r���Z�`
dY3�}�˹�Q�0��  ���]v��C֤�e��m��� �; .�!�R�����O"}��i8/�B%�Q���@��T9]ԕ��|GO���y13�M=�v03��U���uF���\y�
<�E���^��B����I����6y�����z�+���s�D����}		���#T��l�&1�R��n2�KQE�90�K�]|�: �r��T�] G��LHΓy�]w�u�'���@:� ��x��j���8t�5�l�`�kj���4�TE���-��=��Z#��V6&�����/Si�z7��7�y��ζ���ߋ�=���Զy��<������:���s�z�Gԭ���*\k�e��Rq�iK��k����(;�#���K&��sly��[*\y�|��ְ}sm֜�d�/�4g��z�s~d�#) �����%߭5B�l"rMcL��R#����m�M��=���"ok�T?���9(�m� ldC��M�{E������l�o*-�+�� �DY÷j[�<�|���~d��R:�2[(��`����2z:�C�ڒ�j���&�g�o��愺��X.L������՚�$SU��(2`���P�O�-������:ɦ=>�d��e�Y�b�T�5��w����%&c�wy�/�C�C`��ҹ f������d�j�3߹�!�B�j�Z�"��l�$�2���zў� ��&���0im�� ��]e�1{7���{�<��2�ii    IEND�B`�PK   ���X��<�8� � /   images/20128c01-dfdf-4258-b49d-382729dffbb1.png\�T�]�>LJ��� �=�"ҍ0��=tH���tw	ҍ��C����<�￾{-�,X7�}v\׾�ل�*��`��D@@����RG@@]���?�����&���,)����?����p��sF@��x�B�����!�������������lg�lf������"�H��Ky����iK o�Okώ��_�%�gJ$��2�!
��E,M��</'k�P*�LMF��EwÙ�BL� ^������3~~�/���疶a7�j�C �ԥ��?��_b2m��E2�0�R��j�?b�*!~�F��T�+WX��$����a�OF�v���40#3쟇����q�����^��凂R�"�D|�<Vit��x  �H��SY���_22��A��x<>����}U��.���;Q}���!�w�ߜ}D�HZĨ�V,�
Έ��9P�� �j��L���3Q�{v�C�D�ȹ��o~s��F�/������AC�x�IK�hȺ!�<�;��k|	Y��Z��3W�����/`��O�!����឵��Ϛh��g��Mq����)��3��Ł>�A�ۯN�t\

Q(_�@����l}A���E
�_D���	U@~2�T:���9�A�L�	��C��HOx#-��C��HhLצ���w�/���b�Ta_�����e�ɤ���W����v�"��U��& ���5�j5���Gщ��J�gsFtm��}��&��~���n~b��Q���*a���#�혮*?{Ø�;܋"��w�@����=����*2{�� ?�������<��W�z�4������H��hI_��s�����S��tO�q��W�GNc�ot��U�7Ls�Vr0p<���MV������X�t��v�.b�s���7ђƉ���an~a=5���03^UnϽz�*��)��M6����$�� ��-a���T!�=�b���CYGI�u��*@���{�I@>���~yô�[x�W�;��l�?���=*��g�Oy�RM��Ҕ*(�(�⫎�On��u��c@���l%���Mឨ� 9Z��(�f�P�t�+� p����3z�_!�+��a� 6�3�+�O=҅�
�%��1����#�
A�:�Fir�[�P�k���"�%������[�<�����J�[�7r�uՅ�WNݯ����������N��qY6馘�2����B�c��
Fu*M�P%WL��_l���i�����36'�7�C�O2�l!��^�oቔ�W?9�ja8$П��^�?Z\Z���c$�� b���PW�g�C��X{������Q� ZOY��K�糴Z��'v���6մ��2�T�����Uр�.�k�m��-��8���$�6T���8y�׊��M���P�s3���e���Ch��O^��>�`�����)���7�)�h�E~�e��&�x"6(K�N�!oÂ�����������K�≘v}����������9���	kW+���{o���t�ʕF<e,�,��i��=� �e���]�37��ʪ�8P��Q�:X��@��������|I[��{���Ns�w)ؙH�}���C���?f���Ϳ
�*�j1y�{��_r�0��9i� -�o���x#.bGt�&�6u0Y2��N#a���Th!.:�Ν}�ł�QE��?]�r���~>��y6;&B�����)"�^�����{V1a"� +��̯���3�W�n�p�@ �����8�<Ph4]�F���f>���M�)NĭƸ�ۓ�,��4a�5�:���B�@�V����DZ)�%K�EZ�#�ꢐ���2C�2Q"va���hfv�;(��ͬ:�4V��Sl���Q|1Bh��hm�wJ 9 ���GŰ��i�zm�"��^�/�����d7\ͳ�Lѣl�-�]^���n$U(���:^��U�h�#�
|�ޓ�+v�zNr��Dg�M�H��/+P_��j!Fv~>&�D��6� fMjX=e��z�L��I�M,Ԩ�>�߾f�[����[�U�&@B�bw�h7HpO͵��p3I>�=כ�]�T�Eu���8��I�ǳ�����0OKٻ�s�Rs�dIk֩��x�ῥ��ۺ�T�9>�cө4����������AɕX���BV���cjy�I&T�s���F�rU1��pu�77���p�Y���ߟ>�U��k<Y��u���>�!9*�wtM0=g���(0[&���%�#Ǉ���@�~�%�x�� U|��D����t<����7��B��!�ZQ4~4�+���V�`�8��	�e�.UO�c �'�zK_ZRRH@�s�A��r6,�=h�'�<��:���������;�tm�W�[u~G��Ek�=�&�
i� a�"Ɣ�Q�ئ�hH���W����)���٬�����%Z�Q����v�v'�&���i:�|Wyԅ�3(�+R>�eО���<IL�"s���S�e�"��}#Ֆ5�ڻ��]B��Ve��o�"���[� O#�	���
��Qh�I�W!����#�?��r~龍����c�~���QZǱ2An�P*|գ�C�.�Cy��٤ �K���"�:&������.���i5�Q�4�̞����q�s�-��GqY ʉ1xv�j�8}�Q�p��Ò�`q�=���E��C��L��8�}<��&�	A�"&���<��N�郀 ���H��4;b�V@��h�J}��F��1l
$�M���#Z�.M��y+R2r���N�F
��܂w=�Yd���i� �Δ������t-��d��3Υ�5h6	aQ}�A���HF�u����V��!�"./�Fu\��	����S��'L��;K���s����,3��DO+�:�Y��g+�&�5�M �[�^��(SpZ(�x?�*��i{�C�R��������F�� �?�%r8P�q�s�?�**Z�M��B���î�_�`�7�:f@Ծ|�kwk<�����
�`���c���qVǮ��@4u$�̈[F������$8�f+!��bh��#ۘ��:
���v|#��h�C��ô,�Ҡ�C�������V#�	wi�lOѫ���ǠP�|�FO3�pʠ޽�cD���9�䩦9�Y���?K	�7��+�E-�K�����D�˅7�챓�C��p���oj�\F��n������9���#V��[#��W���z)f6�2�G>��X�|Мh�Jڞ}��)OKǌ��\M �-��s3X�U��ՇY#���`�Y�F��X!UMH��:;pN���$�ӄ�X�;�ۭ�?e�[P���dd\�p������P� e&bT������!��Sc��V,i���鷐���)�C����Z��+M�9�9;,�XWE�0�߱�ߊ@	o( �0�8���hu��`� ��������x��S�$H���[~a�-P�'�/b6��_=F�g�d�&I��ٝ˕K�yQM��~%׈��aLN �6un��,�&�0U������BY�>h�T\G�oj\��/v�%����TR��U|9U�7�!�x�b�S���A�y���G���R6�i=�o��i@u���L4+>F�G}���D4��֫#�b��s�`�}8�<�����[���h���^�7�v��
�)RE
!.	�=�<ۍ`�K���>�Z���&=��h�U��<�?$���!3�ۖ�����9�H�+\84R��r�	z�����R����2���?V`�������`�ţ����	�ly1tϓC������߬=aC�2���~�DS����:�c�W`��33 a�l�:��TD[	�	}�a����G�M�.�Ke(s�� ��VZ���4g�"�u,��f氨��nS+Q� 2�)�漛Y�,-��ݤ�Q��\?$mFW������H�����kէ���Ŵ.��j��9ls���?*�tIę��ݡ����"���2AR��-�7��8���g�Er��� ����:��Ac�婦�����b�Q����=*v�a�����9<���s{)���G�pO��uk.� j�r<�\5��*ec6��N7J�k�^��C�������f�l@CB#QI~[	ܐ�N���H��}��r��4�@��#�B�>8d�4�E��v��2/���;h?j~p1�����q�U,� 8��ɽ^���sRSSe��n	��_��Gv�~���2#?�����*9f���#�5"�僟8,����.�7}�Q�"�(� ��X���w�
%?�/~~ؙ6%+?�+���h�F(�NS��H�j=n+�'#�+�z�ٰ~*�6�3�Ջ>U,�atR���$���f��O�h�:X\�����U�'F�1�"'g�n W�L>PY����J�<kx�n�I���~��U��E=�6���HQôe�j��Xy���6�/�i f�7:z�Mc�mɥ���e�������?����G����p��"��qO�\�ȭ6�������s,{L���>5�0��K7P�0r~/���#��_8�Ɯ�@o��nv�I��G�jP��TT,'��<��6K� �Q*�\�qa�EI͖K-b���+O�Hz`����?�ja������;쪹��,>�{��*�
�S����I�ƀ��v���o.ц���&Urb|�a������Y�8�Ug�f"�l�@����͹M�A�}���P5RK�%�^:d��#I<� �zv�W+g��-)+�焥��ba�^�֎]��^��*ĖǺjк,���26�De
�TSչ��>i�	�k�����
�8:.Dq�-�*Z���pUPvmn���3FÖ���KD��
�Me����|h ����+9��.���v��m��(֕�"C��k����x<�,qo�q���P�v԰a��Z��Te�&�6>��u~�VN=��c��+��E��\�BW��@�G!m��*O��*ϛ_�O(s65B&Q��A��r�8 �xj�(\���ia�q0kX.�i�JZ#���m�%�{��������uc��m��C�0�9Gc�k�#m��m_��^�(�vX�p{uH��§)�NK4����FMOƃq��X �nh�҂!��:HB�D�9���u�BF�P���w�~x�j���6�=Ǖ��Q�^H5��Ķ3 .$�����JҰm2l��&X�0e��z:�{"��A�ק�G�'*�RDj�^�PI)����<Q�,y��� ʬ��r���.gU^�ߝM���B�ٱ��J(	���H	��Y~�n�U���n��=~y!�x�X�ᦏ�k���U���/�]��>�$�_�KP\�#��o��V����B���\#�����_�>� ;[�|�u/z&�eM�L���ޘW�%���g����K�u�����(и���R���>�a��:��"�����q�!Zw��O��ڰ�tA�>T(Q���$ēzq�,g,p�4��[���K��C�=�j�&bސd����S�k��+}0`q[��l���W��?/�Ҋxp�J�������_L
�>6�����gj$>!�����J�+fXTC�x�!�m�f���i��~ě�纕ͬ��l�`:b\�����e���ʗoz�o���v�"�rP�k�V,BM������������㑇#Ͼ�^��<P,d������-�H��;�J�����G֧�;���֓��-_E�^Z��O쫶&4@�Rk�n$齆����m���ʅ$i$xlÆ?��:�"��J�z�ޥs���R������Xnk�-gƞ�����E�.4Le��1��p�7�ë��Sɏ?�yh�H�r\��tk12��بbx���4�=O7oՙi[2z�_�sЎ<�b��-��7	޳\����g�1�oߪv���Z�p�ó	-(?�lM?@\���px<���y���89����6��7�x�/�5A�R����W*�&,n�6 V�t��m9��f)�;,ڻ��H�+鶴묃�&H`_e��"��e1�\(�CՋ.����RB݄��P�:�OYw;�~P*�1K9e�n?���s.���X\.�%�FU�2ײ{Wc��,�De�NT>�d̥����EX{kR0���gq$�~�g}YF\-���)��~���'��\�]�Ñ��o�Qf� Mr�#|�])��f��w)aԈH��{�9�:�:^����g9�j�Yl.�ڢ�A�BEΪvg%��k{�f����:��M�iߴ�A��a1��Lx%�KJ&p:G}j����*�n����2�$G:�D�h/�^��Xz��'=�Ş{<�z�ȁa2��'��ɇ>�s��^l�D��ڮ���Y��$��4���-D��cN-��y#Ѧ�7�W�EM���W���� :K�v��d����s<��k
��4��%��
�o<���i���YFݒ �/b&^��Q#x�up��z�$<,�|�4�����e�!�Οr�x�,gɲ|3"������E�,>4�C)O#��]@s�o'��uF�� �"6r�c�:>ۏwP'�e���q����
�`�K��D�؟2��BV���`�w�ڍ����~���L�q�j���M�T�Y}�4���(9�\j3������q�N��/��ļ�-t�;驺�>w`������8�����.C"oB���&6���Y- ��n���͸x�i9�������]����yC��ӭ�K��e�&���8­�
�B���׾�T �}��_~�����^���"tW��i�xǕI�NA���x��m�Cs,-�F�f�ww����	»�5$���q�&�0����/raz(�ޙM�Q�t$�V2��|�L��Q�:���|�V�R��������$Z��b��H�Y�1��s�U�N���E���c�w��Չ�ZL>Z\]���QzW>�<�R�d��b_��/�hp�T�}�zc�M�ut�$�C�������Hn� S0�?J�;zt��^DҞ��y�Z����*�#t�dP~q�a���B�r[-�r&���o��Ufs���C��젃*L5t��E�,�%0#�{dE[�'�)��[���9�ޏ�=�>v��I�ֱáV����/aa(��TRڔ4mUɚi�o���ADa�kwk�$�Аɉ�x'p��,�*0�c[�+��m�咂2?��"?>t�K�!�I"*C�z�����#F|%��!�h"j�s��a]� F�u}j�U���eDu�~���߀�f-׭%�zV��XF��Dݤ�P��]	3�ɜB�:q���C{��`�7�_�lȀ���<a��咆R>4��T4��m��2 �70hͳ������^�Q�c��켕$	�w}�E�dqF!��	���C"�7��쌨��ޢ��� 
��W�;� ���R�kO{�،�(b8�"�����/D<�I�����H��n��l���QO���}c��W�����C8(�����wT-���u�X��҂k��'5�}��:]2m:p�G�8ճ�}BU��[?q��x[�J?ƭ<ZX�+it%����i�8�ݵ/G�o/ʆ�&QT�#:�H�s��x*��&��h�wi�Ň-��4��V�O����R�T=4m�䣐1��7��߿��nS�7�Vc�1wY�J�=q&��-I'�����ya����6Zh��[�}\M*���@f٧N�wl�|-<�KcW�H�q�/�:)�2��!�ǿ��#
7�n^����l�t����khM2~���t�+�a�X塞��}�:v틬�����h�|Y�p`}6�
���G疯��� �t�M�3ƺ�,1�ݫRv��p������To�Jz�������F�������I�|�U�f����7c�ux�ėZ�������r����HN(�Fow�^����i�z@�s,�ߝ���%��x�s�ʓ@�:n]��Z�>��b6VO��U��43�t1Yi��7�?����0���k�쏗B
%�B �7vܔK rx�#Sb�8d$B��C��\Jݐb"M����܁"3a'F�����>/8�.��M���A���H���+Zl+�fE_�k�-5'�{�ˑ�O�Ttr��d�O4���|�r=�}a=١��F��}�1_���H�G��5ڨt���[g�jvzp�H��^{�����[rxLw�1��Л��)��15�b��]/�b_[�ˡ�>�	����VZ���ۣ�"I�Y%��r��q�<_��^��=�X}[�<�=���r9�:լA�b~MC�{��H3�?V���̂�ŷ��+M����k��n�Y�A��-��V��	P҅�O�tM����һ+�%/v��4<�C�ևR�v�l�tߝ	@�;6�y���F��o�U~�\�](��ὀ+)�:�`!��ZAm�,��wfTk��t�I�վ��21͵�Z7�PXK o��� 	�-ɐͯnɘ����8�����0;�d��#֬9��.2 o[-������F��,:��m�B��M��2Hb+�Sra��&�Ҿ	�j7����,g��{79���uoC�b���6h&����|^y�6����|TK�<�%ոc\ѷs`�ه.�rq�����ew�Ձ"�4��XE\�G��2Y�Cfc.XU��	1�q��ּB�Mg�R<X�+;�gq�l�Mi��.?�ic+s"�N1��]"*��j�(��қ]9�J�&���<�t(�ѿ�C���4糖�iY�H�M��8�2Ӑ�����(>��7x�8��slDG�9+.ذD��({��#J7ع��+��A(�e��.�vZž�MZ�9��&v�7`�%�P�4��6��ov�26�\���S���ܟt��T$p� ��nGKpl�

cԑ%�IB�hw'�blSB����*N�S<�L��߀��~�J�����Q%جV�-�F���zYJ��eq�y�{x\�cM�5?�X�廱�����'1�ëڿ��%�zwyĔ6���� k���Wj- Lw3g� Lʪ/�k��o`�s���C���Ǳ��ɿ����Cm.�Sv���l�.�~H.w�t.�w~4�x����5>�YoJ�l���z5
C���g�w��B�s��#���c�蟝_��Y('�����������]U󘡠��%ۈKK��A	�g��6����^�Ջ�ዛI�Xw+��o����Tx8�d)���l�ܝ�as�-�>��ٹ�Ba���#R��V�~�-��B>ɭ+ލ�Z��\T�{}�������0��0�U�u���#x���<�>{�թ� - �ɚ��A:^�F3�t��Լ	0� \I����_8K�J�����G�-���FM��<�c�<����)��=^��*�,�5!�_��*���eF�aߙR����h�]�Ŷ�z�	��ח��f!�'i�����8i�'v�a�t�U��C�.mwl~5����p!K�*ț�M5�9ɥ�p��R������Y�ׁ�	�ݕ�yC`J�%"%I��y��3kGS��j��)�����lޓn�/2 r�FT��Μ��9�LW'B8��##�	��������@��e����:ډݟ�e�� "���m���~��D���>+���*��@Ǖ�������ԭQ���KS���שT���>�"_���I�n֫�ő��E�R�ȚK�I"�k9��%�צܛ(���+$��ʋ��@q�]��G���LA��x!@��@؀�����8RJ�-�(�Zt�f{��%Iр��ݥu������G�AA`��`���2�X��t�5gѡ5;s5}����U�)�.ϑ�a��	�w(�<7:�Zsm���ZT*�(�C�0��9]������h5����7j��)�8����M�^�
�-/L*~tI��pU�#��f�-�
mT�"��_c�uZV}�-�[]�K~�[ݫ+��z:!b��C��%��K���f���O��Hk�YG5�F-/Gȧ�kN����#��z&��p�m;\|�q���;��55v?sW� �ԯ�;H��+7��.Ԝ�,�y��ݧ{�؎�}~����yG�\PH���gu҃^o�����ྸ5N0�����>�<r�ú��$Ֆ�;H���G�Y����w����ȸl�^� ��=�0���N�'��Y`zЋ�a��uY��)�ͷ�9:�{�5�]�O�U�{pbI��j���� ��5Hx����΍mX�<fg��o�����#�����qU��<�V�E�.��=��By�t��1I��h�&-&*I|DK-e��d��c���N�7Hf�;~�V�,.�n�p/_v�����g(���e�Ge��(�E�ȗ0�+�:���s`LO�����!�V�i�E��ט�����p����'g�m��0�ٲ��
�~k)��!i�,σ䤤 ���т%	�G�J�"�i��*u���=��sJ���p��Q�&Jj���k���?ܤޚ]z�l
k�v��J��{�]��[����a����B������]�Ǽ�_�&Iel�b��-���!��^�ע�?�o��)]2 v���X������㝗��g6�|5��	�pw���B-:cW������4|{�8��XxԶkZ�u��ZK;UԮ�Ɋnsd��,�R���·��-��P���ޡ�hy�XU�jP��px�{u|�y��Z#x�,�,�l�{���N�=�#�\�Ì�B�+�@*��6�$��^�������9�4C���c��V�;w-�2'�i>���L���Yk�������;��{��o�}��"b}�٪8?����X�g!� �K�A���q0[Q�gI�]���/�ٴ,��F��M�]�Yk��Z�q����?�aMɎp���M�wr���9��15��ݰ����ڡ�(g|�������x���4�5�H����a!�����ns�Y����?����ď��R5'Q�#a;Ơ'�/�8���ּG��`��=:�y
�l1��յЬ�8.��Yn�� TBu}�y��	�� a�mW��'�*�i�|��&TF7 �D>��fsZ=:z��x W��>9�p���:�gU�'40¶��b܎�3P�{,�R��>�.YW��K5땻?��3����r�y��{�F�XZqA�_�����ϓŘRLA �|���t{W�Fyh��"��R:��)9��j���\F	x�{n�41ƒ��t�>�}Q�<~m>N����-众n�ݺ�L�>��۶�4򺻖�"���Z_���r{^�(iL�e�Ğ�@~2O)�#���#�y��]g���K�IAT�QqP���^B�������:��kF��Z29��Q[y)�s8 Ij�����G̭��HD7�?.5�p;)`�~��ב�B����2b$".�R$�G�����̓�W�V
�Y���O���K������"�@��3�moв�
u7�AHB8H"9=;#���Cr>P�lR'/|�C��OEW�V���x0;�Z �;��T�L��5g��"�	���br�w�-a�QT��M����cr�6،L��@���t�ܳBz�G$�u�7.�x��ǡg��R	�8ۛ�Q�L�(Ă�U~N���U��v�4M��Cɾ�V���O0��߷'R~�[�O+9Ob�PJ�oղz�V�k�ѫ��Vz�=���V����b�geܟ�QK�T���VH:\*�MA�Z�a>>��Y�@�}8���2��hS�l�P�,5߽�p$�\���na魰�-�M�[���)��N�D�t��5z��7�oIY�,����l�6���lbz�Vo��O��i�E��I��ED��W����G��Ѯ�>�_���L�:�	�,M��6��eux���f��(���Z�%$�h��A|��tJ�o�P̓LW� `�RK��y/���ƕۉ��y-��6r��G�f�%��L�Sg�=v��P$40W�@�7TT13sP�h��\C�j�\�Kځh�g��f!��ǷgŒ��߂�������4�vo���������b'9jkgCm}=<Y�'�N��Oi	��d�ŋS;Mrb�?�_k�D��� 3��������~8F�������ִ*�|�q�Ǉ`���8�K,҇���b�68�5���>�4(!�{���?��4���Ls���HP����lG�m_�@3�W��H�{�h?e9��{�2�
&C;�E�	��>#�I�ka�0".���]��<��ז5�٤�I'��q�#��:��q�~��,��z.�� 
H��
{����`��A��7�ZI�P���@C�N��a�ՈŴ���N�����t?�)c���%ZS�R�D����}��j<&�=Y�0�K�~�Si�lY젅z�Ԝ��fk���TT�qT,�
��?�\�,��s����%H����gwS!ok,��z�>LP����V{Qcm��/�]0��[ào�$��+��X���Z�(ӄ�R���3�s���/�n�FyD�a��n��ޯˏj&���v�Og�Į��_p�+S���U��w���Ǌ*�e6Yj=�;{����� �)�%�jd��c"����_2��mF���&� �*m$��Q�*�#y�����r�z�]zO|D
�%|��?(@�t�(��j����8�<UUwf窞�m96�p��� "F����+�r�jQ��Z�^m�e��x�Va���ӭgx&2�/����类Y�SO��9��:��p1iP�ֱ��`ye4����b(۹��ZN�/BJ�=�"zws��8@q����0�A�d`�<��	��/h�-��|h�
ӗRW0�y>�[q�����ď����d
��Tv�9]�P��>�~�I�G����\������^c�?M���7��n_���	��K�h�2�����w��~=�Xc����=1��♮�����.��a/��e����[�K�����\����-���d��/zy�=�R3���k�<	����t2�A�:��n�]cT�q!���W<��JF��N.J��t��m�]�Ƅ,��|M����ĵ��Z�Ϟ�Yc+9Ǘ	B�NR�ve���{Z`����h �ٮv�����xJc�4yKc��_��Rs��өQ%:-���Β�����y��k�:��G����#����1�8vCK�3j�G:��ꮮe�3$���C��F��f�vәf9v�����ڷ����p�S>�A^a*��d��'�+��X�F+��Lܜ	`4�M�{��o�	C}4��=J�m����0�������uo#tKt>�S�e�o���g7a����n�oSI�,�&��9��;��P���Wh��rB��*7D�dB���5���*X�G#:�^,��M>��<�f?��X���3-�	\}�#�݇aR�ݵ���b�\�X����~�y�lϦ�ͩ�r���F1d'��H#Z��x�q\���TJ��Z�U#s.'��!ޠ� ��I��q�]�x��j���B2����;a����6}���Qկ3�\p�6�<�d���I6����M�{ڰt��ɑ::��;Q[1�;��Za=�mE@U��Qs�����c�q�E���`q����� *�V]�Gm�'���E~��z�L���K(j`��z'���#S���إ��p�|�Q��O>(��b���k�F��z<P�z\�g-:�nU5!"(@-�kv�2�I�P�x�����t��]$��{	}Z:J�pO��2�Δ�A�~m��R1�AM���tE��K�S�y��h��Uƀ5'||�� %;sچw?�[�o���ΜNk��������J� ��n��P���[v�����}tW2��k-��3�)��0M�j����_mk�,9��"��4y����_#��X<�Ɔ'�TS�@��"�S�wJ��7D0����j�lk�/��n�x2�T�:��	D%,n�8b���]F-�M����10���e���w�I�[��*N�:�=�[��ꚺJ5��̧W��y�z����mJ�Q��N�&�&_�r�4��ѦQ�G�iZ��[B�D�7Y�B<vrSO��3Ӯ�n�J������*Y���jQ#��F���U��abb��|�Y�26Ė�N+Cmp�RL���w�F�@)o�W2�ϗ^�r�	OE�k�MI��S<L�K��y|��������6#��������a ��c�Fǁb
��O�jw:|?�b�&�_�F��+�=
ro'���_���[fښ��/P56[|����Ʋ^�����5+����9���� �Z9�q�����m��cD4ð���!����q��󰓭����ٽ~{&�z3-mK=(Gi�f4+�߀A)�O�X�*ϥ��`-�2��;VaҘ\�?��xq���<Zڭw��wy������s�r\M�9���dl+�'���O�i�V�~5.�|M)~��=�~_:w��dMk�Qx쥋������!$��I�o�j�$b��Nm������h�V��:p2�ݩQ�u�,�UgP�!-'N`3}�Oθc�(++�]������{�V������U�5]�bG�<\Q�ծ�(��@H�&�+1|b�h��*7/�B;����C�w*R[��+���p�Hz���IIk��k�_�ܿ��i�N=�\J���֌?#�.D�4d���#���܃�S�Χ�E��޲Q{�QݺX)�)�ǃ*�4W��yמ*���4��C��O)u���$���R�����+Iع�y����� �8���V�5Q%=n�;�}�>􁄼
�0�:2E�~7�K����m������6H�-{DL�;�t�X�COݞ�O�e}��a������f�ǌEf6�����q�beY��*������.���d.��aX�S��eA�Kвh����J/�A��ۜI8�>�DZʩ5�ksv�R���F^Dm�Vg�����1O�K�1��ȍ�L/�A��_������ʻv%J 
��r�E�.]k���.V5C~�4��B�@�̖����3�=��X<��ǫ���5��A͜;�E���;�!��:���"Y�u?��8?��EJX����K������ٜ�FS���1��j�����W�o	2��(��~yW����U�B\d��!����"_������͟�哫K"���]���7ΐ��ǋ��x'����֞��O��d�F�|�̣~_�T=MvQx�@XH��0a[ɉђs�e�9��EJ���T�
r�ʬ�u:|�x���^�&�ɪ�ߖ����&���w������󩍕��UШ��W3Vo!0TGk�gJ�j��@��9�P���s�0�Hūӥ���wh�szhw}&00�K\��;�����ǝMŤ~21��}��1��}�����E����Q�P�IL�^�S����%��'�Ȥ�>��VM�0A�}ܷ[]��{M[<�)\��Y/�=㸂:�����oC~��|H��F(kx�	|�W�{��x�麻�S���?���j�Dw�6�ɐ��R�$]7�%�������cC��Gs���� ~�hQ[�>����֟;I�iƔ�����ȯ�kI�(���mU�����w�������?*-	�#vf���<�8�@��W��-Xd�u� �65^�
ܴ 5X��j�������v䮧͜iZ3"��8h_>
I<ƈiYdXF`[��F�<v�}�Le�)������4X�n�co�.��B���-v�;9�M�.J���� �`�8V&�y��9�4���Ǧ��$��R�S���jd�L]Q��2����Dj�c"e��� �5"+�#o�d�J���N�j������Пf��f����6�����#xĚ��y�6Rә�|�6��P�F��oȞ
YY+7�1�h��� x���f{8���&�(���W�	ܔ2��4����ܶr�i}����ҙ�)}O�QZ�R10Ojw��!@Ǫ�ũ):��*9�N���5khrt]N�7Z�|k��t^��\E�qE\�U ��x���&y�+��n����܇9/�5�����M�ae�U����%�u�9�����z�/��cQRf|�B�=����8�+|��О�+2�5��S�4|��g��#�Y��$�F6���6�v�:���#��].f�j��t�>���لTzI�:e�]���4d{]&����Q�˅h���ȓ�܆&�A��㧁��P������\~�J\�7��|T�����Ň�8#D��_��k������L��3Έ�h �UJr�Wھ�;f^{��.�ly�����E�0�����Qf��v�@3�<��+�n�hA<5xP���۽���cM-h��B���h�ɋ^kɎp�WGN2�B�r.p���D .�n-L�y۬���&C>������D�#8,W��M}fv�(uj��>g�DZ!�sgH%0tV>��Cj/�LkRE�W��Z��o^�A6)��#2_��3L������P[�6�r���Yi���&�j2�{Ut�٬ԟlsw�u\Dȹ�S9W2����0��^��ގF�>R�N��sA�����u_�+8)���a��ƴ��r�/9H�#~������p�\O�-#���͈��\�C��D���#���'.�5�)$���M<���윚^b���ѫ�"$��/�,q���'y?$΢+�Y�h#K���h�� .���{����-���i�g���������I�琷_�X�L��#gR��5!v�_ӫ��C�VViO���O^�6��~��t�����o���}��92�����i�7R��OR{Y-6וw�z�+:�%�v�p �ߖ�A�
hΚ?t~�d�8;�@��Ȫ�3I4���f!�ԁ��є+���t�ʴ2Ē�Yv~����z밪�/Z����Q������HJJ7H��H须���q����}߽�_>x�^k�1�c���ݾ���E+�����D\,�hY�	�y�7�I�d�q��1��jo��}��ܰiW���EX#�vP���K�!���?͍Ձj{¾	�:���^����ncw{����n���]���� c	��2����NYs]w�w��T��@��Г�	�\�U�c�n O��������ےRKxX�1F�Ø�S��C8�s�2%��ܕ��`d̖*��р��$��bd��>�(6�Q:r��Z���b�k�qXiF�$`���<�ǆ���:*�f6C-�
WFh�Gl�yl�q�[W���yu}e ��A��.��m��/�ڝ��F�[�G�k���5���ȘO�@4������+���p!apC�� a�a�Gr%��a���b���K�=�,�q��p+�a�L���o./r�T�p�CC�M�q��m#����Y��UL�|0%V YR���f��r�ZfP�^��M[vZGn��WQy����]�;U`{l��ڈ/�m�'��c�MH5Y��^� d3��`��8��oI3S�˙��:v�#l��L�#�'.�QiuY+�]�C�bo[�y. ��;�ӳ��-��u*��c�}Sse�£�ao-MY'���T� �����V�yn4+���F���ntkK=�2���d��{
�{���fBl� ���0����0�n�ATe����e��)9�~����Ŏ��7����9~��INQ8�*��x �������z=O5�~�s�[�v����ܡC�`�LԣC���faw��e�i��d�?���ey;�	�y]�ᶻ7�a���=@P�;��aM*z�1��{���<o��{e���WtA�xzO�/<:��FXB��ז��J��>d�
q)�Tl�q+[�����`��d��$Ԭ\^�
���q�A��!�޻t;=�p��kN�v���|�X��
�B!�+*_Yc��b��a��'�E~��,s�a�/�i�k�ͪɌa0�x.଻M<[�'h\���(�J�M����R\�N|����4��V����ڔ�x�P�~gfP@}�n���̈́��|�g�!�F��G�'��ZPU��`���/	D�?Kl��7�G�]�O�2�_F�(�(��]V�k�-�xlC`Kb�r���v�|}�I�>�7��	�zכ��h����<�l�\��j�'3"J�dOiE*�J�\b�g,���O���'�5.v�@�y?ٜ3�kZ渹	��!�l���]o��w�o�1�C�� cr)"<�yI8�S�ڧ9�&�m�(�;�`�%�����[v���*{�r��nc�)��v%V��{�[&���Pe_G*���g�p3%�i��v䑅�m%t��yB�>D�.��!Y��B�B�Ψ"��Y�
������e4��X,-ϟ��Rvފg�����:������v8�/;�)���͍i��#Ӻ���|�[�pd=G���V��#r����37X��ٞh����E��ȕ,���AO��ޒ�Ia��=�+��)~w��4�ϋ0�n�L�RR���ș��K�^�b�s�G �)s���dԝ�aP��E8qL;�aM�
&��s ��(��yS:��'Mx�,CY�������K�Hag�0\!�	\r[M���r,]�O��)�)��4dd���N�b\ l��B���<I��Rİ<Q�a��ވg�D��;5x�)�f����p��(�DBm���Fź�:��'��V���S��X�~3o�,��=�'��������Y1��m�.iFW�km�tR~���;N̦
\�x
s��j�^�w�<�v�u�9�����C/#�>+8v�9���ǛE��%Vlli�3�)����b-Jǁ́����g�iuY\k�%�Ȅ��%�m�����AI,'��삎ʎѳ���w'�\�Âu[>����%@$+��G��!ĺP�rA�LFt�����U5*\�����:z���8PH�^�[�m�A�,m:���@S�G�֧ߔ]���á�]n����=�Y"->O+.6����2f��� 5������D��7��)���!�ե�H�oo\��M,/k�j>r7�7Z�dh��{�?Y+���9V�YN��ơ$��z2��q����x�F��>�Yj\8uA�^uZ��$%��6y:���}�^	h:�L�+�M�~vl��?2�D�ş:��8^'�K���'(���<-����dH[��f��X��^�=ۜ��̚�3�ⴵ�7� ES�5��u,�|�+-�188���m��X�{����N(#_d[33���B3�fxiV<��C�g�,�����>�I��+����B�ׄ�5���-�_���q�'zrp�bcmT����EmH�~��0�Q�ɼ�&9�#�j����| ;���56�4���K<>��/�40J���/T��z�'�Ƶ���-����_X-ػ�\��v�J�&�ҖTY,���\��=�z�IJ�x�GD}�
�1�-btKj��m�����N!ͽ�O%��N*�[�a:`�.������A�;s�gd�6er��{���T���=�D�$��Z���c�9ʭ��,�ڴ��NFbW������4�i���G{�U�O��0�U[K��N�b>}���"�>lCL� ���[f3$Tm
A�^�R8ŤeI5,�����<m� ��+{M��lb�֔<�-
��a)ƍ���Je�����л8[�;im�:J�����f�5e䎚\��l�[�7m�b7<��CW�	�ebf�!�2��
u�44�}p�^y���*���n�Q�)Ѥ��PB�P�r������)TςC�����w���m�f�F.r��x����a��A�So*Vzo��}Z;���V[�Ţ"�?�'N���Z�E���Gs�,�|���Q�ӫH�*�z���A�H����7��1�Ֆ��Y��=���}�pd���o�7�Ob�j�������,
�8ԙ��<��.�{p�T�`$�m��H	)�o����[��O�tD�Ǯ�7��f��w<�<�{ k!ģB��_^$�|�����j�Hd>��� ��3d��i+�͘��|�f�C��-���Jx6E�P)��9���n���F/#��?�D�S��{Y�．}��ꩼ�]�듥����{�D��s�F�#-0���ٟ����, �^ f_Y�?j�S�&�\:�z�Oj�����Տ�0�\d�"�&�����Fl�<e�W�fF^���v�g�$�0�D�)�y��n������g�){���\��s��W.{g=��$U�:��`�u!���a[��2��&\�'4un���:pg{����[�M臹�!����{볰 9����b
��t&�iՔ�}5��Œ�m|O��k��mH�er c"±A�^V���Fȃ�W�"��k+k���e�Y�c/9�r�)pw��|S�v8�:��@����C" �^OM�!�Kk�L�\:m޻�*��݂��`}�)���ק���$�x���\,/�Or�P��r��Zk�8�?������(P�
�U�������\����#"���23�hב���.1��bKM)�p�i5͆{����V�Y���N�J4��>�3~J���C����J�������7�[}!��/O�ԒÍn�5�k�hmE� ���|����3�p"���LZw�,��o�#�$���jY3��o)���<r�2J�Y	�u���g���/y���d�8�H]3MeF�,�D &�P�~T1�R�Tm�F�K�~�nC~���H��`�^�K�����qi&"W�s��ঁ6_O�.������Y�O�r��׈��H0�9���Ϗ� �^�=�Pr�X�L�7G0���D'P)�z�1�F��LV�w�m��|0;��I�}��L����|�#�^7�yzL����<�H���l��/��'��-�n%��Wz���Vx��Oi�7-B���Q�����в��kw\�KS���<��+�d�s9X�fP�J��]��G:��n�Jؠ;K���B/H�Rc�T��4w{kKI�`��Fz���U����D�B�zC^�T�����x�l�`@!a�R?1���F�r�&��=fC�ˆ�b��������	��q3(@k3�EMZ���ߞ�V���w�7��wD�L�n�KH�y�:���Y�/k�>Ӂ����0E�S��_KYPUw�%�a�)�7?����3kH���mn��#���>uh7����`W)��ꚜks���w �q��Ed>�	:�����g�;P�Ȥ��I�7�p?�	����+C/���3_���c�/����t��q�%L�m��>�)t�3v$J]����|�1��4���x�����)��l�Ib�Op�l:��_�J�Gx��g��<����c���uԝ�zV��44�,��}���7�0Bh��B� ��2��7j�O.@�ǖ<a��x�����eyQ���yң�^�t�Z���)�?t�p�S����`���|�P�^{O7���c��nA|+Nr���s3��� {�kP���w��Oc$�3*A@"����!��kX*� ~�a�3]1��y>��]uS��K��>6�DG�H�H�jف�����I���h/�M<`c�
�9�E�%:Πb�a����,B�L/�+�R��~v4�!\�Z�,�Y���o�
M~q{�)W���{�q��l���pX��^��u��'��� $�q��R��q[�'�2�C&k��x�9��������D.��&��+�v,���~"e��L}s�Ӳ�=��ZXqw��n��i��E�8I'�e0�a����C��W���:n����`�w;�������Hv{t:��]L�e��n��GK����K���������㓘��:ewݭi2��<����r�!u�t9�s?�ov.Z��V�J�a��.,���ޟ���쿲�:���sW���~�S��I���GR�/w�<~��5Z2��%��aNC:�^��x���^�%�����A���Q�Q�ʦ���*��ǂ/���F �v�����?�����������_Z��r%�*��*4�N��tMܢ�x#��
>O�X��zfF�o�reY���QZ
�0�QE��a���t}g+��vK���+|E�y�_�:��,N���c'�'�F�D�d\�Sf<�ai�5��B���`e	C��U3�מoԥ�Ҍ��v���B�n@+�GJ<�/�]敿�խՋ�ף9wͯ����Q�)'#/l� �����Gw�TW^I�b�M@e^'z���?��u�@5���gq3#�9������xa@Q���耄,�BL&���b��̒To�𣸖�5l^.m�0_S/�}��0�ͺ�Ro�YJ_��@��4x�źP�ec�����H�R����V���qi$?�d�L�*5�z��[�Q<aB^91��L�e�A�r��N��Ը'{����a��U�^R������E��`1�H���ϳ�x��n}�1EJG�[��;P,��K=DՔ�~�?H���s���[���K>*p��J�{o���4O���IR�}��d�a>Q&��4�k�x��G���[5a�]�b���}�a��ڣnow.�p�1=���g'U��f��<��N�l��]�-���!t���I
o�"��nWk�Xԭ�>_��a	c��o�����ޡ�V{׳݌�:m��t)0�+�ގ���L�5z���D
�_�)�|�r�'����{Ѯ����.�^�\ޞdn��1���v�����`�ʭ�_�"�Op�X�������kMز%�g��!�C����洴38��U��9�&[��0�M[�SG$��y���k'��+��쥙���!�>6%�����y�Xţff\��?o<
��~��i��sTn�l�_&�>�.��0��A�kw����;3�_֎6��/S���p��r��J�i�T*ٞ�0.�q�K�8�Oj~��&�7� kR�24.��.H�V��y�lK%4�e9�O��z���Ǹ�w�=��px��j�k�(�U��+�S��3sZ�8{�>��0����C�_�����y��um|����R���6��5�/A���~��0	�7�F�Y�&^�b'+HO�ӥq1�je."T��E>q�e#o�1v�`�����3��N���I�-�kCQ �]~�<%�:�6��%4�t��#�����8���K��]�A��ΰ(��#[������ٚ<���[�.�m����WP�Cߘa��&���vɧߏk�ָ[�fD9Ò݈�b����"YD�*Z-E�>�[�y���Z�`!~cB;�e���h�I?��o6��:����3��S�`*s1���PX�я�(#�̨y�'
�Lbr��C}��k���z��y��P�/F�e�"��RL�_"<���{�<H��Sj�	՜7d��X���!A�*#����9��Cd��
��[����a!��u������Ma�*�*������J3�,XS��
�Y+�$]ߧ]lNNe涑���<^lQ^A���}���	��^^+~��:�|k�P=��DO�	���!p5ɾ�R�H�����6PF5m;v_������m)�0��~��1N�*����Z/�c�3��aI)�S���О��~;i���3n�o�dq���.P����0�6l�ًI��	����u�C���YO Ē��r8.��HA�w������2G�ss��l��׺a�������XG��Mn���q1�N#�M��𴏮G��r���=�����_G[�W_&yQ7/���[3��H�C"s�"���Z��a��>Z�Ѐ�;��?�C�(,+ښ���Y���H�DMI���h�D����Àj�xм_'Η��c����e�*
r�y~Z�w8�'"�SټF�I�h�����%/���Cp�3Q��F���1�
��~��a�|շ(g�F�6K=W��?�LM9���(���+z�)!�0�F?WU?��%�0U���9�<���#m����+��4�3:k�0?�5�谋lo���4�73؟+�W"��Tş+��<� ��4�c�.r�[�]���ks8EM:c!T��h4���B0�'� JT�4�.��I#KqL�&�	�G�xa�ը��C<�#�X8k�3�#�麚���Hös�'�����u��/7��5d觲A���z%�T��>�3:BYՍߕ��L��Jeւ$}�K�+����J@��j��$	a�ʽْo(O}S�Io�q�(�+h��IPe�� ���K�FF����w,����tUn��/,ve��8J}�\�!��VRI��|�~��O�)�}_tkr>!�`.�E�cV>�DWN_����/�?*+�
e� R��.�n]HX6� �ؔ�\�F@$�Á|���>m�kA�x�.�;L?>���h�7�i,�i���qCv���v�r�O��\������ϛi�!����t�|�
i�ʌ@�}��;�?�KC�e�Uq"4���r����j_��&K|�y���>��D��g[w��@��Q�^h�,t�����q�v^{]�Ο�rW��]�J��L���L�����:_�g�����V�'��B�� �<�K)\�)��M뗏B����ѯ
l��a�i�������Љ^a�`�ņk}B�;�S��L*eIjJ9�죉�N$��<�-��}5�J���$�^;��u�g�l�-{\��������Q��l��-�#��+9�Ro/ڀ�9*�tC��Z�FALs�[��798̅����^r�3K5��l��D��*l<�D���"���|������w��d%��Sg"�s
��YeIl4��3���t�ތ��Ļ)�glF���9q�4�i�*�-wl�5WjO �x�A���v�fH�YY�؃�^��	GM�c^��u�Z3�"�.���`�̂9Qf�ж�Ux�.d�-\��˻B�,SH���倇�ζJ;b_�c�&}.��6'_Im�¿��yg�tT$�͘w%�ꔾ��f�FIF"�J��a=���>�|���E\PՑ�Q�d"Vk�v����a����bdFX�	1A�|[C�NU�Y9g�o��u`�OU
F�#!r�A���+���Ϭ�nת�'��E�M�C����,�OE��6�dքB���q���P��p�gbo�C���fD�hζ��ǵ| l�@-(����oI�a�)�+N�h����J�G�+�~�G�h�8�Qx'y��&���26���ߏ�4�5Ʊb�i��&�N�g��4�0�b������汍أ�����r�g�S�mc�˻։���1��`+_�|��� $J�灞��-�b�(U!_O޽�^Fr.���NO��(�̖w�13�_}�Yk�P)έ�J�4�7��pt��*Zݎ;��̣~Ji��O|/�U��Q8�-��?�F��j!q:��*|�Ձ�X[���uu���<XqK��5v�x������I;ƻ��H7�7�N�eX����dx�r���~̅'��N�R��'��#�.���:�]��d�jэ��:���z*�(�T�zsNp���O�Ք�3ᙡ�
W�J�>'��l(����@�7�㖕����@M+h��ʴuT}4vs��NX�g���ӝ��{�p&����8!ҫ������Ę��`�_ÿ�o������_���w9C���kS��w�#��a+�7Ͽu���*��T~�utO��Z��X�EC3ʸI�N^P�5 g�M��Zb;É�*��S�l�m!v�`z$J�3uۣ���~c�3\fwJsξ�$��Bu��G��l�]Dn $!՜u`
���i�*S	��e����B9��0�׋"���#s�M' ��ۭ�o��ٝ Um�	�|���c���d�+M�>u(S�d�Ǩ�^���c��h�I��	0$�rF��!��l�6S����_��\�.dVmH�d��aޗ/lE���2�=��j8���o]����(;�B��+3=G#��?1�JU]��������~#�{Qx�f�2�����m�OI��Ҹ>�@���7���<j���uh��L�*t��u��*f!I'����=�_����H�V�Z�]u��H��)�];�������T�{����v��������yv���B6y��`����Ap�ӢwHmw=�$�
��h�''�(Vca����Y�m	�t
�Mfrg1a�~��:ٗ~�j��%����7g9�;F�k���_����rB.0��- ���%�}ɮD}�Q���R��X�CJ_Zx&�l`�T�h�T�ݭ������&�{"��Lܥ�	a��	T?��2ί�����I��@GO���,	���0�e�Pګ�-�,yiI� �j��^'>��_Ӏ�4N���CC��<6qW��'����U))wy�����)*�xr�;�@J' ��b�'k��/��j�a��(��A��wnn�^��fw�9����9�qx'ָ���	�o�"����gGC����:�ϐ��+@����ȑ�f���u-�Y�9��/��a�d_x����lV3�<Ջj�VR^��^&�p���� V��s�����{����su��h�a�7{b�����(5=�}m�'�~�+���`�FׂF=?쑄��U?��?��c�%�֗�k'q��D���-�߳%��+��?�N�bu����֋ "�g��
we�i7����n�ᴖ����)���@�<Ϯ}�z��یg�e�Ҟ���C������0�>��]z%a_<���m�ſ���ԩ	M����}��*���\�wG�=�Q\�I��ma��d�1 ��l-;	
�QA��z�����~��c�ےE�\7<�j�m(��+1j������3#Z�߈����+�����3+v�+�����̐d}���
�}q������A�8_4��Ԓ�V�����h�y���g��� �r��;3ǼF$����tP��7������MУ��U�VV��Gû�A�"8���k l`�^T��Äb̩ۃv��c ��1��|Źz��, ]�-O�eg�Y�����r�ݫiW0�wؔ�-����Գ�6����;'��&Lb��1E�(����٢G�0�]��'�~�?����,�ɼJ��2�dTU�ʽ(����U���H��)?�X�4�8N���h��g=��3ƣ ��Wˌ���z�V�TيO�*�,�M.|������ ��!+�z�`�,�h>��)d�����l�QJ=]P�2��4�+[���8��{�r����j�Q�"�h�`�U�Xtx��6�KvX؉_��M�=�-�\�~˗�nML��,S��(�pɻ�/1�B�G�z�Qն{�{^hAy�c�$o�4����V��x����LlJq���Wm�`(������l������nw}�aZO��L\�>"�*���ÂB����|�`�A��<{*��G��G��%*��LU�P*���y����N	���1�9qMb�d���;l�؝s}d���X�c�ޡ}�����A�uZ��?;�{7�3k ��LH��*O>��&FY��j�xM�����K=[�j��b��G���جʋ�J�pN�j���n��g��f�lw}t��ʦ��|Q,ժi�`���.vF��~5|x�G2���T��H���.]������� }Z�(N*Wʅ�/�oᩤ�I�F���~kL]���	��.Bm��5�u��A��@|�����l��������df�N1��+?r���~s+���@�X`/���4g8�UvbgqI��/a=�#z��	K\��GiŻ�|�㽋�Z? �|$�H>װ�� v^q��nT 98�$Q��
�3Q�
��wX|�����c����wi��S�óy@�B��:*ꪡ�w���7�_@(�慎+a�B�3?
�������i��-<���_9�<���|օl���B]�v�D������ɿ���A�[]:A[�v`�}��=��.������馵�pظS������἞�͟����%�TṈʿ�t�F�DԲ���ȓ_��,U�]�󀂮�����X�24:��k��� C�0nI�I�0�w�;�#K�5�k�~��6�HS5����o�������1�I窶�lm<�ʋ����q
ҿ$�T��v�˫�6>Z�i��EWHI��.jZ���o��x 3"����g��>���_��C��;�J�R*.'��i/�$�~�Vw
;R�;���I����i�c���sVe�`7���r�}���-�G ц�����1��i#� �amQߢ�EqP�ĂdX0I�YP�_���Wք_49���t��[��|��t�1�Uu���Z"��U;S) ��=LR��k#Ӯ�Wϖ>ܞ�Se���+Z'�����;|�-�������w�΄�V��7)��IV�D"�[�}��۠���W�C?1��9��%�$H�6����n��g��ɛo�J��FJ����3Y�d9��#o��Ԧ��M<h���_F\B��Ų�����8��]�m�w�h�]�:Q��`cK�:�Gsi]Z:]���V&��]_��V�T���J6���KmԢlȤ���s�ep��yL�B��T��� ?_�+��1�c�z4�������L���?��&��@
R�q�P�h�����Kp�H�:��h3A�a���s� ���@>�}Ac�a4wH�����U0�s!�[Z�q�u��R'y�q���ȓY��v&!q&��*\��P�MҲD����R��p>e;������I�)�9�Ǯ���^��6G�lhF�Q���{���m�`)L�@ݜꥯ��{��=�Zw�t�LNa�gl�n,�q\���5���Wz��0���Q�eե�XR��:�á1,�6��f�ʵ�f�+Nh�_0L/���z��̏j �����Y2���z���P4�wL붓8J�=��d|K�&���<p�g}c3~O�p鉳���}r�5er�v�|��X�Gd�(Zq�Z{����z��z���uI�'hҫ\'P�V��$�^�g?1#^�M�4#˺LVSe}��Vp�_�'�����@��q�w2�	������'ǐ��D�{��3�B���桪��A����o�W�u}�x"Z����#�t�$��)�*�r���ę�S�	��v�qv��>Nv�#뜄� FNR�����Ϳ6�6b�,�5veY�N�sL `��L����K��I�s<����R*M��K��	=�9c7����Z�=B��a����!�͍���b�=����r����w��z�_���Sj��	�~��j!�����cc�Q�3p��XA��K�3�1�7#4����]DL/��H������`�L�2`�z,��LB�m>�X_�y�X��F�z@��-:��)�~�^J6옛]�_�GE"�X��E��?S��7��v�st(�����KWe��j��(�%63W�ΐS�X��}F�����u;_) ֽ�K|r�L [�|U��hk�~�9���a��b��@�_hb>>l/�5�4�GE�5�˙�ՠ`��πE�#C0���x��־$$��pJ�R1�$��!�Q#�Y��m}x�����6�JBހ���P��ו�L�\ `����)�dYYM��T�C+ҹ��ӧ�H!q���g�0*յhT0	��z��^��^-�S�(� �x�*赆^��(�������7���1?)r��7��n�����ak-��#	�d����6����/�ӻ1v�_�mpN��(�*�U?�pCey�-IT�n��#SK�����}��@6�'cլ_�B(V(��ú`~�"��.{2�?�����,�2�z��G�2-VL@�^�[���-����CJ�X];�$%�<�J����r'($B
�y�w~�˙C�P��L���d ��|�}Vy�+��vM�6�RE9`jh#��{��3�����,\�O  T`��f<�`���~@gVQ���U2�s4@y�� l1��WP���~j��\�mB}
8h0��Z�%/u	%��o3&�9)�v q�T\P�,[�o�+g���E8��,�܎�T��������;�w]4�J�ߪ��'�u7}ͧ�Px��8�Y �׸�Q9�u{���lU���9Sb�R,H��O�Q��:�q�"�W'?��7�
M�c$Xn\�'̃��/+��%G��5��Ka��)DCt��Qv�y�:u�Q�ڹ���JU���yI�A��QY���*
�@�y١�˥�	µ�Wt��?�;ݘkW�^������Ϳ�9��eGI\�H2(-�%t$�dqIo	Ȅ:�f��{���%�iq��X�qP�	�<��9�~�N��W�R��b�fz�}{��RM�"
 pq?��^ų[SY-;��w��,���0@�|��oTϐ�9=�G�kQ�Ҍ�z4�U!��1K�?�<��G���-�c��T� = �)8���p�d�&��8�-7p��1EG���f���zǸr!�'��'��|��*iL9��nT��+꿒���5_}�bTrx�>���-�_8�~֡��.�sf(��au��"��>�H�����I�����KZ�����P�O��U�F<=¯B�~2�u\$��s����\���N.���Sxռ��5�s]c�7_�	d�'�IZ�6��kÃŗ�E�n��ru�)9{�DF��@�a辟?�X���'�Nb��8y8׼��( ��W3����R��nC����<`Ja��_V�z03���T��{��bҁ���|�%zA��ՠ���ҟ�"�Z*������e�ŹuSղ~Z���e��Ū�Z ��ٳ����P���v;���,���������Jz��MT**��ֵ7���c&�X�:}�"��F���P�� m�/T�����7Tl&�S���w�*�gS��uvv��-�g�,@�4�� 28�x- ��%>������?6�Y�L��7��� 6��=e>�5�0cI�9��#V|;��cWಳs�"Ω�K�G�ë�ڿ��?��I$�w�a�<P������hLO\��`X�6qv&��K{!&��^����gM��_�ELx��(��e�1��[�.��s��rc��yB�tz��,����t���u*.Ux@��U�g��6�m��@�"���R�BR�7����{���2K��a�����E���P@k�����`�</ʌ��j�y�y��&,|��ֵ�S���8M���U�n��T��۰�9~}� u�/�$)@"^^�+��X��.�YB:�F�u�<P����?�K�^�VK>J[w�Ki�FR)����P����xc¿�� �$@��g�4��{�V���F�g�
�f�^�چB<�f�·�Z!Mer
�A�N0^�άR��ﺞ�]�c"~�����g̫�'��T��u"{��h�g"MQE��wS��J{[�Y+���7���̵��&���o5��>��y���R�J_�E����-?킭$d�: ;���9B���\h�s���$`��ܑ���f|=sLI�l��E�'/�7X���C]S��� ~�0���e䯫�&�b'y�s���<��Aj�
v=�X�mWЛʺ��/-�̠���(SB��r�g��o���N�|�DU+V��%1DL1>��G�j��i@��r����~ZR���Y�@�;+ZG�ӳUy"(���	۔ON#��F�w4Ou%� ��JqbD�cg[KEn�â��=���ꄷVV����(�|R�{ǲG��Y_>EX�!!��3=
�27S�E]����=�VNH�Okhԝud8���!p-��lG9G��¤���u�%�ǀ>�{���v�}�G�fҽ�	��w^�j���#��B�0�k�KOv($���S��� Q��xK���d𘊇��M=�3�٦Q��r�|����i����X��ي����OKr�̑��� M���\fy�l�I���u�/�'J�Y�a���ԟ���H\����y�E�6�)�W(�~�8VP���`��(���k��d&���V�P?�~�^/��~��X%��׈����Ue0dx/��S�e��+#2R�9���)�}W�P���!т�"ԉ;����Z���P�C���h��:�����ph�=�ae|��|�	���pRQ�P0n(�kݟ�ҥ��K+�ۇ�4�t@k�U�@~�[E��FGrU#�:N1��Sk����j�FT=_���=iJ`�9�l{���U���ɗ3�1�u�#T����Gj�� �4�B���\b��B��؊SJ��Σ4y8�	�w�=1��E9���3���
I,����Xv��W�)cǻ��!�h�I�[����3�-i�~���'�ϳ��bgT!��2�VV�"�=���0C����r��.�ɵ�n�!u�D`��ȃ:6�^h$�-hb�p�#e��,�sC_H۰�11)�.��K>�6��c�q��˺�Ͱ���d� tʴ�SV
�=��73w�Z�o�s��@� i� >�զ���Z�^�(�N�m�`�Pؕ0N2��1��e�Sdg�!�N ���d)��A�e��K�����i�8#��zݿ�mw���xmٖ{��?N���ݑg(���pG����]Շ+�R(���M�x_c����^e��^8�9m���Ԥ����
N�g��4b�z��-�}$�����δ�aK
�\�d�E���n��v�xZn(Ը-n.d��Iz�"�oP�3/����w*��ǰ�n��\�� _�%����j���+�/R�$	$n�Æ���̻(�z�xF��a������vZ���0� -��a��6�P��Ox�:��"��:�Г;H�z�[q&��w���>Q^�C�+��:�7�3p|��|���<�G��Z���Xd�����j���������CL�����}T������Ѻ�R+��q�K�&Xp`g*��2����t����s�Oj6<�|~��=�g�T�k�My���`<͹H򐽊5{�>�J�6(��F;�9;��O@_��R��8��i3%y���i�y���h��|1�-$o�:%"�Hei�sTh6���*Js�QkO7��`ӓ�rϐy��Cx3J4��7&��yLX�θ��?M<^�+L�j9�'��zqw���|���C�#x�$��td��T
��� �	����Wv��u]k)�ib<��By����c�ky�������>����F��UrE�@��C��"��8�u�Pլ��A1��(o�ET��'�o���GʝS]��[��\,����>�
)�Q���S���"�V��c�S����a����Ƀ�)���á��6,�M�?|(?r�}:¸$Y0H�b�-c��a
����W������8����R�r�����N@�r�/[t<���;�+=:��r��Ɗ�Ejl1h�eR�Q�l�?����
���f�c���ae%�vS�o�|m?�v�J\a ���H�J��GF��*Umǻi�栞���o� �j�,:b�iÏ)��}���S�l<*4n�*$��\�i��OghX�4Үy�~��T�4 �%xd���KE���h��gHm�l�g���O8޾v� V<G�Ύ�)V+}Rp�D|���&����F�
\��$���� g�l95"-�ٸ4J>9gDَk��rs�u��Uтv�4��|ѕ9|@Q-=�t�F��	w|l��$nL����P�:�Њ���"�=��-�����0����H�������"�u�<߬��I��!����P#.���~�+�v����Kv�P\�|��*���=o}���4���9 )�Km���5��iO&�Q),�Ӊ�\��zn*���.H�\��˛Xf𚢟0J�
ß����Q�Q�oS%�r��x���h��$�'�R<�y$/�ɘ|�u��'I�|�E}LR5�ꅙi�Kk� �imj��8����I�������qQ6�ۀ�ҡ���tw,!���ݝKw	�%Jwww,!)ݹt-�t7��|�ߟ����3�\1s�!��nG;����0�F!�+�r��Y44G<�tm+���&�A�δ8f<;��%����c;U�r��F��=��ݹg蚙�a�P�,�إvnk0rϨ۾�T�e���z�v��wr״�n��r��+������g%AT�aQ��/3�M:oS�بJ��?�%�\��^a5�
�	>���>ȼW�jhy:~��a8��W��F��Oӭ��Z��9�I� =H�o?J?�'�ޤ��d^�8pm �c������_De�᜞��(,��6�plkftk��?Y�i���Kq���!5
6+�FʈV������+ֻ��Wz��N�4h�W�������)"��@�4�����K8��lє�z��?�L���"ÿEO�8p���7Vz(J�������"��ϋ�5>�S�F*�,�6l9�o }Z�t��UN��mmJc�U��zr�ƴ �Yr~n1h-��ټ�@�]F�Yui��"D޵[�k&�ꨓ:w�	d�=R��5��x��;|־t���z��i���{W��Jed�����9��"���u1&<���ӭ���9����n]`�	j�Hf��ٚ��z�y��7�C��hu�~\%���Q�5��W~��5^����"͕�s>$���B���/�=w��_�˰�h�"�FX�`|Ap}�r���fQI3����5��]_V���l�"�g���۰�!d]��)B��~����M8�y�K���.�0f	�<2����;�lp�5bB�����U��������Wb�1��_�.�˪�C)���z:R��q?� �#��zI'�f�{ѧ^mŦ�͍R�4[���X�jKcvy���ʗ��N���߱��i1���m���G���`�᝔t8���zjt��0(U2���Մ
u�8����߶y�8E��~��I|���-f�j�5���La�$��Z���PÝi���,�3yۛ%Ko#lD�,B�e�Cw؉�M *Z��yC;�M����4y���E������	a w�z��:��� �+4��!R���b�e	c�+�א~�1!��_���u��z�?�T�&��*����K�dZM&X2%p#�c�#E�	\�TP,�]��ŝ�X��=�5X4��@�I�TZ�2�X��~<%t�笨)ƿ� +&N��
t��^[�p�q}8*Ec*�c?Ы�!�ʪ7tr3�^�+:R���\�>J��b3d��ܰ���. �cn���:�K�_Ƒ�>ke�t �y�A7G�S2���M�BC�$��|!W�G���P��Y��~���*	���pl�tEE���VQ��'��W�7	>E�_�d��������B3�yA����|��J����^:���x}7�����9�\�P鬠a��[?�[� ����{k������(�=����צ��5����V`4t�����>�d�#a����8��|�!NLEV��P)�I=���i�UL\Q
��nfң']ϫ)(B\88R�c2Q��^�!_��˖y�����y�i�ԏE�HR����A���ho�5���@o�`fw���ͺ�Y�oSGl��V���lI���.zu`2W�,��fŒ�i�
l�����@������M#i)��������"�w:v���煻fW�O>ElG�����j^ޥ�x�k+�.�٨�Թ�A��^(�뾒�zGY1�N���i:;��uネ�ƥ���B�f���S���n��d29���y)��DB�$�D2�����ؤ�5+���0FR��>{C	V��a�77��ٴ��CS�t;\�xĩz� �{� )x�)t{Q&a �y�z*zYV��_:6����*)�/.ud�H�TaM	�)�ғ҄�TZs�+A�F6n�F#z��N:f?�PY4�ɠG���4���_�'���j�+Sy�@�2��V<�H���y܉DԢ��w ���Ò�Cv&c����\X��}��]Ɉ������S�.]H�I�R�o�٘8���I�u/Q����Dǌ�1��b�>�@�ױ����c3����~#ǟPs
Ƃ�0�*�^@����A	KO����t��=��/ű��XF�ݼt԰�@�MeV8*�����O���5�2�tC��n�V��f!-o��Q��s����ɠz�y���ۈ�l���h��0�lG��4� �x�'����Y*��S��e�JS��LI�~�̕6ԧ|�ܷ9�N=���(0��⋭�6��d*��.6��4�|x����k��}��s��7�{�Q� ;����$���.����r"�~���OP���T���4�!�X�n��ˎm��h*��4웓|Ђ�j
Pb�����27�ؖL{��y%� �NL�7���L����m<l̗Z= ѡ�~�ʘS��R�G|��|�|���}�C	󾻁��Oԯz2�*"\��yu98�C���?C�*U�F|�o^yN�	-�R>뻨�(4��?̗����6ן�]ZV�P�z�E%�~Ǌjj��B�� 
�i��Sŕ?�i�k;cB�2!�,eԑ��ͬV e{[zY��������cGA�b@#��M����b�����g羆��?E�����eS���<K	Ѓ�
��<��G!Dm�D/P���U*s���$��2�OpY�$/�ǜ=���-<s��k:{ùe���7b�n�W\=T-��O�y�D�Y���5"ٗh�@�*i�mS+�n/��������8ep����.�k������q'D���iW��A��!~.̽G;`�HH��R=����i2	=��woߏaa����%����~��q����eٝ�m$��P�fD8�]0��� ox9/��ۯ�^�Nޑ��Q0࣐_���hr��=<�>7�ih�b�X�֣�l-�ʣ��� w�\��v�m��7Jjr�O:pн3��"��L-yS�K+���4�������lA_;o���X�Ijn=-��C㛿+l�sn�p�U���E����I���),�Y�s�8N)WG����h8H<��sR\4� �U���M��]�?Y��9���ܶH�>��A��`�2�Q�^y�nF_p�z��v����og\���7�s����d<�;2���A�����\���;@��Saz`��AT��vGX��%���~s1$��s��<�}~�N`����rx"X'B1Ѫ�+m�}�PoM�e[[��%�j���5[���,jڡz���K�
��,+�Ύi#yK�r�.�h��$aq����t�;�t�p�t�Q�9b�\���A��?�u����e�����&����e#
��}G�?KL���mi2u�>geຮ�l�_��'G#��A�I�����]�,��!2��"!�m��w��=$�ńa���Q��o}/ྨ�����G��z��Wz�>���y�:mߌ�s�����mƓ6���w�{���C,S��	
���o�Q�6��2�rZ|���cOe���UK�DU����Hc4ݧ��E���>Ͷ�'�b�e�Ԃp;۰W���y��0HOЪ|�G�z���&��{f^��I�)O�[�^6�l��3���h�e{���K'Y��Wj)�k��?���K��������H���mO��Z�=�ܑ�l����>��۸����})ë�z��nL؏Q�W�;�Vq<FIy��D3ɹ��]�-_!,J�)K{�X����X��LYC9�<ar��>�#�L�B}����N:��cv�����q�+�J���-9�������5��/�CB2U��#���i�sB�*���7KG�3މ ��t�[��[pa
��in��s"T�ڶ�yKd�׉0b���yn�kkz�����u�]hՅ��u[���*�gO��|��t�^v���+�ݱ1��I��yx�w�Q�vHZ�f�E{�՝�S���֍΂�Ya�Vp������0��p�oF��u_��|j�wy}�P����n�C�}�Lb����v�R�`�i���Po����`X��I�Ma����j��AN�/`�~񑔵���@Z5�Ph�qw @hnh��*�6�J�k/�O�4�k3#3"��aģ��ї"²q����M�x�H����"�* uy���$,C{:�$7���kD{)⌜�-,=|[͋W�Gb�-?T�+�݀�-&��m!����*��ow|q'yJv:���;M�i��B�J���Oن�i��za@�>�,U���դ4��T?r���ֵ�[i�*�pv�L�M��a-b�\���40�ka^�"S2/�\�Qn�#Okw溘]���%-���	���Rt�9�h����Q J�5�:ϼO^zP�i���r�V����	fn�p(ؓ]�u�����U*�[��������Lֱx�Y!�)�ꄯ����a��оʏֶ~�|���-k��QrM-��5jPH�����R�pD��U�`݈��������@����l�50郄-I%�#]D�-Lqpͭ���>/Z�^�MmA���LY?�5��X�sj���g����3��t�_&C��lӊd��6��8߿X�17��w"J���������p��e-�&��&;0{%��Ӟu ��&%/��eVC#���L��P�+�;�����?��1
�L]�y£U�C�ì,=�68�_���Ȳ@7��.�}��ѕ>$u�Y_ʹ.��P��G�j��~���rޑ���Ew��88q�#�����"�� �+FH����(7�,�_8����"l�_���|\&�
�1ȣq�KwR�����]1�RȲ��#O��K#�y�Uو���Ǉњ.d���V[���z�~x�z��ښ��Y���b��P�i�ƝB���`�{�Ȫ�%��E��vA
Rf�NX�w�4D�����w����P,>���W�B�_Cawڗ:}{YE�X[���9�]�x�攂H.2���{ڌ�g�[��;+�,">"L�^4�tG�xަ�V�t�h44ܥ�ϧ7.9���Q�<E���;Q4� c鱒�x�GXn8W1�'%� t��>��;yFi6��y�ni���$)�haA��Nߗ��i��	����Б�ǍϝX�p��jG3#���i{"^D��gy�;��f�~�N ȝ�`�8����nSLIժݼ�9\��LǼS�d��l"6�g���89�G��/�E_m{���M�'��w�RY��m���v&��Q�_�BoQoTv@W�Lkߍ
[�Y�&Xj��Pi�7�.跕}�L�/3A���}-d�z�}�Z�X&�E��<��gN:)���V2��lxh]�QP*�Ty�[�夤������Þy�kV����#������0���� �&�xD�|�kˤ�wu�� 
�hy�)�[����`��uX���E���C=�L|��9�o��t�{yf^�TH���0�������I��7�Ǵq]G�)kۢ���F]������-���a�8�y��a�S�{��'fͷ�[�GC����ę�!S9�p�nd&m/D�*F7/	v�L��/|�p=J3r�;yt�E L�i�ԏ*zK�<���5,��j�'7P}�Ł�Y�u��T�b�Ɇy�]!A�|^��J��2��O-ao���N��\��$���d��{
�6k|�EҢ�țû�@x����)q�/p��~��]^v� �f��L��mx�<X֝r`���,�//�|���:�%�Xj+���������;Q�Y��Y���Ol4��0�:y���oG�)1m��9���#h��_�������~iꪏ����2u�G[C�ՠ��;��������s\���(�Msܪ7��C��ٚbNRs�!���Qg���j�x�4'�v�Ԃ]X��{sƘle���a@͓4�~kQ�hꋘ���������B�g+$�+�������Q�"1L���ؙ\���K��A�����I����rdRF!�O�"���q����J� ��dP�y�K�F(la�!7 �3k���L��Υ�j����j?��ᔩ���2�_Hƃ�|f�AD���U-�Kz��[e�'���+��L�h�GJ��=��\�����*�KV���/o���7Md�g~4Y^�G��c bj㣘�^���F�#����ԉ;	됗9�ۥ��<:7O�;�-���עUr�%s���3���T�l`���ApԎߍ�l�����)�a���5~��c_E�n��|�r��Vm�\_�Ҟ΍ӂ�))!l��r��&�Tu��#�'vFU?(w��;�f��In3}���;C���t�>�����9Ԝy��y���:|kr=�,���J��ߜ�=[W��T����[#�@�ұ���6��fyL��q����Ve_�1��r��R(�4�'�n�m�z�$�v�̵�o6���������Q���G[�at��Ӎ�v�����	s{5j8��eJ���MN,�i�	�h�K��0Zps?��G��J9H����W�v�l?�q�F�%��Fcӣ�J�Ci�(��l��/���5}�s��F�ԚI83�9pD����,�T�R�']�`.c�V_��=Qƞ��nʥ/��J/b��|J�!E"J�#����dD�t�J�~�����?�<���s)n�	�X&���Zo��TKzvŸ�qlm}sV�f��VdF��ZZIG���6��k��Po\z3�4��Q�}��Z)UD1
���I����{��o�u�*v
;���5֏5܍n��[�~��r
�T�jX�lE��)�\�L��lH���&�$�vC���>����.:Ѯ�%��i�*1<��x���M婹�{g�0p(G���>"���-�g'�\Dc}��/���]��+�6 ��:w;_��v3V�#S>�P������,Sq��y'�Gǡ��G�����5LU�G!w!f�=#?2�ŭ{h��;\B'�%���� ��@��H�����(����`Ɔ��֏M��o��ǚZ0�af�������ibf>��5�x��og�#by|��ǰQH�Q����˟�1����\R����D���l+  �@��ͨ�y�I�پQ��x��3ب~;)�9��H`)��hi޹&��� ��K󮸋NX_k)J�n���+x������*�誎�Ք��{/����Y@������J��:�s��a���R�t�5�m����'�t���ܹ�|�Q	s��w-ٝF�{v23�κo�d�nQP&nj�ֲ�$��Tۚ�"H.6��؏�|�ƭ�pch��'�D�l���g���K�s���0�[@��v\�:�!7��?;��m%{O���;-i�h'{��}"�Q#����?� 8Hذ��BEG'a�A!֚��.z|��>P�c��}��A���ݟQ�q(���9HO*��'.��P9�*�)`

ͩI� d�
�A�x0��ڑ��@��D�}nY5���Y0)r����l��m*і_5he �LD�ɬg`{�v_�S��`��i����&Ri/�<�3V=��Σ}�b=�ؚ-;W!6B��B�M/�y�F�Hȱ�]%�������2k��y���ת�ΫUb\s�դ����T�![;�xD��:�p˂��>p�ћ3]�r?��/{����y���$_����&G��5��DO��_v�a��u�z3R�g�Ht�+>g�R�4��
��z�� �6Av��6������M�E7:�Z��#q�屦
Ї��2�5P�!,�hT[:���29��y�� ��g�x�co~�4yf�z�3[��nT����R�$3t3�1�鬧��u��N�@1Hp�$��,�/�:17�D��J�)���s�*�͍�"�2�p3�
�ԳO�U_��p�g��QՆ��y">�<�;�2�@�ĂO�'�:a@�İm��_@?}r�˴���Y<��b��:*t%���ΥK��y�o��q8
0�Z�M4ŕ����ع�K�۬¬y�k2��j'�w��J�L���| ��l�Z��� �����{���Q�M�����E��ף���rй�0]�dUߥ��ジ��i�b�ۧiV[�ܣdB��'=��e�5�Gj��F�&�.b�1hЎ�\i{�(Q=Fd�{@?AV���n.z0���ޖ��:��DJ5�����
���#Z]67òp�Kt��v�E����e�LΓ�����/�ʉ�mM5Ko�Sp��ɲ��l��Έd����b5N��W��r�>���:�S�3)g��b��7jsĶ�dۉ�:�>��BI.uK}z����(�
�w �w��D��D��XzA��0'�Oq�{�+�֑ʘ�����uk`�}
���wfB��{R���R�50|�J��WI��cR�ҽ���BK�#p	4������?Z�$X�����P�e�lG��IJOe��VQ�ܫY�KRyb}�����K��1������1��:kp�R�(��R��?lu�R��|�vx@=}�� ��L���c�b�B������?_��ׂ�R��yè�<���f��1Y�5��A0@Z!�8�8��z�*�4�n��7�����b�$�w�f`��P�=Nތ�#|K~�dq�5-+f����o_Zh͕C4x�>x«��hb�����as��S���m�*��ž��Y�A���_�o�(sp�S�y��=��S��<9�= C]�"���*���^�QbŢ{-YP�HOǟ��O�細|"(�a�2\���6�LC�����7SlS��B�ӻ�oܝm��(4y�2|0bpڻ�C���� E��0QN�9��j�ٟr$�5ؽ��dLd!��a��2�
B��(�Ff(�0es��
	��ڿ&���.�Z��c�������'I��[���������p@	�l�>��@e��vO�1oHǇ�"f������s��~�ό�h���M�`W7u� K@5������nYmN�H�"M+���_`9jq�K��;:U�e�E�n&>7p��Ri�:w�em���&�ڇ�^����[���yw���A.a�'*,N�o4x���Y�q���Qq�1�U��yU;������.�u�93j��@�i-�W���'������[���'�tfF�Rݛ��/���uu��k����<�R������m8q��'��ͥ�9��D�#��A��D��Fǁ�����Fn���k^���&�5��8����*�(卦�7�uz�+��z��caB�Ƶ q�Q��6S��G�����_s�&��T�P`p�6"�K0ѹ]�Ź�0��d�c�`��)b L�(ڂOcE���=_H���B�U���՚�]}�}�T��+��,�;�
����TT��i����ϼ(��N0�9��Q�fj�� )M���\��d� ��O�u��T,��B,&�or9�k������T*��D�m�#p�b�⡵�� ��?�>�������MO~���U�z�T�5����T��P��1��ض�}�ov�B���_&'5W��Qǎf<�TAD�ԉ�Ɣ����� 8�ݴ#X��<ƈ�i ב��}��b7(�c���>����e`�"����x��y�S.�J3��!�ЫN��k�2�i���q�}�$��}p#H���E�sWtPE�-�]���"�=Kh���~�����!̢.����x�f�%ͮ�#?e�b|�}��r),�����:}tkw|3#ؑE���xm��2p��p@�[C;�R��fR��n��xKu��)X��퓙w��Է��EAn~�`�qL�$�ƪaWdN{?#@���L��.u%WǕ��iV%u��=��ez�����g]_�l@�lP�<��2����e�H�pyT*J^
��:V�z�I3>�4^������X�!�ǿQխB
��,ˁM5	ۅ����
�_A��Gf��ڙmJ
7wZ�rS2� ;1�7���3��0�?y6!W����u@�vx�÷!�E��d�0��H^Q�_���Aӫ�X�)k��A��K��=A���t�z,v@�E�-�~��~�����H�f��S?3�$�v��#vGR�HU8ga�'���1�X������BN��U�݃�
��(q&�[�v��-��-VYj���ǧn��7��s��6�H9�y��9�A��4椄8���~�/�@���[�D��9.��1��7r	_#�ȚU"G1�Bxٿt:��^�2��Q�v�M�OK4�9�˲X���]��"9��%����vU�]o3�|�w41�.^��'�ǡdvv(_$���Ӱf�|1)s�@��0��R������p��P$���]DW��K��	�$��{^���<���;��/I����#s�=h�/�4.��lY���ާ]�S���Q#�5��X.�ǃ��y$�2YQCm���3#U\�A�5����ڻ�Ng�.�zyv��E�T�|U��c"����f��R�y�r`�O��좉7-%3K��Vh$q�U�{$Hc�c�zm����K����eÃ��7^�YVL<׫�%a�w���M��+���RW�Kw�`��V�\-r7vq�t<o/`q|x8�����Q��A���/D��2��~���+�"������R��;�p�h��gm�~Y涵-,�kt v�?U,�>��,o�P9ma�����˔Z_73�p�:=��ّbD����J��8�*D�e�*'�,a��|��i�� Z��qp�*�yp��H��/x݀�(� �ܧ��y��{T�����Ļl/OU���~�R�hX�z�c�{)��0�/Ȃ�T��l7���_�Q�v�w�[�(��a��;jj��Ѹ����7|}9|�V<����7!���WMD����m��3E������;V:p}8O� �� ��u���o�B�@0dl��_G�H�3�aJ�Z&������t0�:V\��Yg��&l��t�C���N�zu'�
oD?�-�����*i��ҷI���
f��q~M؜�I�F}{x�����Q)���S���	���錣z�@W����Җ�O|�i�adQ�f� �Ҫ:�E���7���g���T��[/�m��t��4&�l,��b��(�m����섷�@K��atY�Ȃ�nI�>�dls���+-IuK��W����?w��P��+D��6р�=L��D�kA�4&�P�5�#���_�e����д���5b��J<�V�c�k�ϸ�=R�K�1�o��d1�|Y�����w��t���-j~s#-F��Gi@���C�`V+��y}�
�Vz�ymD.4m����u�ҷ��"�o��X���䛭W��k4��#��)c��GuO/�w��]������u��� �Ȼԛ��]�O?ʗt�����q<����b�c�v�ǹ�/���z��z&!�i��q<�D@.�,��Ԭ�&�%̬'E��<�� yp�^b��m�x���������h�Y�R��_�I��M'�n��ŁN���@��ڊ�]�լ��-]�Я,}mXW]?��x�n��U��fl{bg7�*
x�.��N��*������PꎸrtNg��5�\��wL}^+��n�`f\y��s���<�>����6ΤDrR-c�=���#]�)�Z�zX,�_c�
prf�*&ic�x=tR���w+�s�*�VG�9uq�5�TY��?yZ��(�{	o�JL�YS/e��hC��j��Q�H��g�Õ���ao�PV���1$U����55�Ln�ܓ��0jD|��4tp�4U����>wp��N�&�:ۀ�:�6ȅ�P�;��ǹ���n�e����Dǭ��z��Х�yQ������4'�������}�v;[���xV�d�o�s6V�����<�Ljb{M4A�즑��zr��������A�)"�`|�1����X��h�T�m��0e��=�v�ZMEyN0"��ʿҾ��Ni(,�@ 2e%��%h�qX��[<X��XQ�'B*���_�7�p�`qLG8(6��g��>�ؘ|�(�����m������XUۨm�"�V��
�5p��� 9�}��r����p#�����5ߥ��6�r�Vm�BP�����*�b�$�h<�O�sq3δ�`�� �x�b�ew��r�)�g�-n7�њ�����P7)�|�q%��/Դb�a�8��·f�������)�X����aa�S����gkLɎ�fN!L��ZQλ�H��e��_wz<ig+�|�ȑ�و�q�ஓ�ڌФ�;���:i�t�P��cdG�-�r���S��a�{]���Üe%��긶���&�/(ƽ]VA5_W��r�`q��e.Zk)ܮ�R@M;���/�9��[Q��Y^rm[�R���d�O�b�@K��m�=�kCvq��ϙl~ĳ�Wn��c`~ת�Q�to4z[{
 @}!����7�GD�:��w޷c��+Go�����_�G��a�M�~V��=��K	�cC�\^�*\$�g��_�؁J+xlt��%O�*u]U���
OcP2��C�6�Gg�YM�
�1U^��cT[�nd��Pj��t�:3"L\nN���N��2s0�������d�,$G���c��p�<��1��Cu�S��Mߓ�ia������BtX�>%K�r�H8��8��PAʓxo�~D69����͍����֜�.oW;��S
���
�]~��uMX8)ռ��NMqE��+�'?�e��s0JZs���P�z���v���A�$�o��t{��46�ތq7VO��7�I7��4�t���33.\3��_�U׬����m��Ŷ	O�|�X�kX��tM(��|qo�������ᄸ-3a���u��������9�����'�a�Lҡt���G�@�����*�"R�e�iੜ�n��P`�o��@Fٳ��n5�Gi�D���e����'TR!��z���S�ͪ�Q���2�Y�'	ְ���g[�zu|����g���w���m�n6k�}s�^P!��ݒ���;��1i���^v��C#��|;S����O!wz�.�c08	 ?=�J�A���T ?�.z U�צ��⿞-��n	�UF�aɪ[��2���8Eh��9�93Qњ-��kuf-�MU_OE�σ�e�P7dl�8��$I�{x�����:)�R�Ck>N��F��^R��Z��n�t�`�w_T��Og��L5�S����9��cߨ��c�\��]���OZ^s�?D��]���^���]yy�#�1ލ~XV���U+�(�Y�Vi�_�֡�Y)�fϸ-f~�:�s�1����B�f����H�5Ȃ���f�\+���A�C8|�!sܯ7�4oRo�?�6M�c��1:�t�F�o�	ʞ��G�;mYŬ��Ԣ�B
(�AD7�Km/y1aaϡ����2��\��>�l�V���m��G�;��q�ޗ�*L�Ynp*[:��]�뀱n_�~�!7R��	��Rc��۫ bc)냘�Y~����)��&���d��He�[u𖄮��s��P������[$ 4�� :t��Z����"jQ���H*�>8�n��(���D�kdI&�hlEgň�C�k �B�3��������W0�� �*<��LA��Г��o˾h$�
t?�芋_���
B�=Ïʑ�j}�ȝ�r%���:\Gn��&#��1��[��!��ђ�t]:Xn���J+[�����[��h���v�_�ݼ1��s�U������:J���%�D��)��%��e�m`Ė��f�o��K���g�J�zvvA�S�r���(�Mߛ��.��}��F�L�u�#��3�:��k!o&g������d0b�es.� 5��N��&�z����;&�6��+�n�Fr$i�i�E9*��"��P�[+z᧲��k�A�R+�%="���SH&��C�	��>yz�q���a>h��]�я!+�u��K �k82y��zTy	����������9��	�/���Bp;��&����ā~����V�6�A.�W��r��z/��Rk/��v���MJcp������ǿQ1�}��w��iϰ��?3�C�'ܦ�Tx�4����}4�z�[�c�����n�R�R��N��*�W�4Ao����=�%�� x��>�Vc�pg��m�םB�@��X��7Ε슊��U�f���
X�����Y��xH�^�D6gN��O�m����P��S!�@ݯ�O��l0]���ֺo��W��VދƟ������3�[�O;To���l�szX���]��Po稏��v�~ѶC��.�h�g�;��:fz;��$�z��Ӭ\��?���ul��r����sw��^�׫&�����a�A;�%W\0�
��w�����ȥuh IQL�t �V���o��b����.�x$��=aG���л�=��$'݆be���jV�Ps'������-7u�]E�aE;T��B��rjP|'���X�@�;/ۚ�o$��������Wo0�;���Dr=m�~#�����J4 _4�S���D/�Z8�?k��in0)<+��7���M+��3�}$�b���uM���^�|\�ͯ��#�{<���d2���T�p����42��8+{�h�R���-_���	��]��͵t��
�N�6������Ɍ#;����!��K��ۇ��R����$.��{/������eܼ����ȫ+]P�~U7�r�z��A�k롯+�ׄ�$˲��_���3-B�������z��gi�Ww�-�������#��ɿ�탽���}Ж_Ǆ�Se:<����M0ƞ��2$ջ>��oFL�1���K	H�����E�ٕn��T-�҄B��=Ĝ0
־���a��h3q�F0W���'(힝�y�G�ɍ��/���#�>E��������������;ÀoK����0B�VWR�M��G�qD��?[�ԍ�Q�(8k�K�J��&LU�u���3
��&���%_���׆�\oؓ�0�#Td��:W^6Ez..����4 w0�E����y��T��b"�!/��sr(m����?��V���ÒٞnWŤV�-�'A��#��\Ϋ�5I�<���[�o&[f�߾F]�������x J�/�B&�P��e_Ƅ��\ă�ߪZ�v�I<����=r@������87ܺ�Q���&�
��ؙ1��.%������-�W��y`}�M��cu�/�WV���5"�\4i��������UZ�����ʴa�����n�?�N�?������l�R%�T��#�J[��o�ۏSa�$��6O��2l^
��^;��Vh�T\��q�E�O��|��f�Mz�i���_���ykqt0��Q�$�T�Ӥ�#w��M@�y?/�����������a6"���^(4*��Nw~tD����%��IX�ns���J׶�u� 7f���Sa���Q>�1Al�W��X]�sE���ey5��*͜<e�̓��H}�N3K��i������h5cN��I��&M�S�5wn��(��e�w��~R�[��,�໡GU�͝����(���,���xH��N0/�eOWr+|a!] ~a	1
c���M�~P��`����Y�ӟ�j�.�2ŭJ7_،�����K?����V&�VY,�N���5�w��1��v���z�?'����꼵F�A�.q��Z,Oi��&Kd��)F�����.`c����{4����sGt����H��W���-fB���i� ���45�pPd,v�����g�f����o���l6_�&��.O|=��ȓK��)d�H�B���y��4�{:"Ux�g�7� �����Zb���"�i�c�
�ų��v��sМ�*mB5hv#x�<H�A�X�<d�)C��5m���|��h&U����>ؠb�I���p˽���p!�ɓ���Ҫ��$LЄZ�ytڅ����S#��Y���Y�5]~s���Y{�p^��̋��N���\�^)ܐ����S
Oj��K)t(�%]��/�$e�y�	��Ų��&g�%�����>.�sZ��������;�+�@z�8�+1k�o��Q����#�����]�|`tC16%�fo��j0��\��r*f�إl�I���C��b^y��.a�e�״�(27�ђT����c�d��=�7�/Cc��w�����WQ/�У�铅��%�9�̧N<Lr��UD���$�B�?˚�h�i�e&	�U�&�V�_�'�ۭ��Rp\�d�S)?�=���f����}>݇���rk���pA�S�}9�pO@p�E�6���9rFw�����!�H-����Z1%�%Q�q'̚E��VWDǙ(��'���SN�p.z��k�̻]��	@�������r���/�ǂ[~:`a�W����?�}���Ω��+cgY3W�������~��ֽ���%�8��[R�/<LrF{x䥲*��%*��E>~��U�e3�L�ܪX1������}��� 8����1R�����_K�@���Ylb������nRa����V�\a���jd�3g������x��o�u����V5�t)��g��yZ!Mn7⢮������B�i��Ԅ/�n����I�_�I`��ߎ�U()����M���磛�䞛X'��,�Za�F�֔,e�6�Nb9[0��dA��[�ϑ?�%B�Fe�a3,%��h�y�M��רyC�V[�>���,�q���J֕O���1���1b�{։S"����*3���)A��@�Sm�i���Y:l�x��'do����*���ɺ�_my��W"6>h��ҵ���`c����uTT��7:��"�����JHC�twwww�"�����)5t%�������}��޻~w=k=k�?�Y��������z��{�3���|�����+(e^�{�4��U�=�2Z�{ l�'o�Ux#el��`b�����:[�8��蔸?�{ jI|\bխ��_ж<��t�@������j�V�$blm���2)[�a��њ4S1w����Q��+7za��Fn��<���^ث����N�D�@�i�r�'U�b*t�+������E,���[5T҅xu���������}-?$=��5b�g��.nz�G��3t%GV4��C剦t3��I[��¬kj��%�}�7���Կ�B���o���r㈪���rg
�'�'婞�eW�owW��s�$7�������>���y z��T/ x�%���'��T�u���6	��%p5���?�(^v�D3Y��G00��EZ��r���a�Q�`W��%�A3���;��1н�� ����W#f%���i"�7h����'];E�74>����Xeph��_v$������N�̝��є���q"6�@�9�R0:�I��f�v@E YU�u��nXm����M
�י�+���iEK�A	i�h�?��`?J���"ޢ�le�w�5���l�`8U~����U��U+�����,�w �������'zɑ08�D��qM����.�j����S*v��>z�?�{���}j���T�W��G��V�0売�Eq٤�$�7m���-�<�4���{sQ�D�s� H��`!�����.�>�P8U��Q)�����և�/����H�Y˧9�����{�At;�hC��?1y$s?dx*�������4B������(^ � FrD-�Q�|/Q�G�o]隷�5�N�*pnǞL��nB^H�b��r��G2�~R��(ds�0��05"]�>�D�Ë��r���,<��Ro�}�5��V�t�0�g�Z�O�m)���#���Vd���]�ݴΙ�$��=��ukݥ�k��ItW}��R%�ݪNz{���x+V�	G{%�����W���������K
���/�뿠�?�����k�yJ��MR+��.��'\`���I�\9X�,��胊������K_gS�K������`缙O�QA���� �b�&�Ww`���;�����2��)��U����>3W���&D�\���B����Z��4�?������/���o:�z�ï�����A���Co5�,֋9���$��L~ڿݵ �1�����@	܉%�#F�q��+罉����A���>+?���$��M����r^X�Æ�r|�VU#���S�}+e��O� �ZWk�z��$����D?a�u�����kWr#�i�2�j#@��=�A������	�D̨�}���AG�=�����F���%���'5"A����P�}�m�]z˪�5W+��Φ�5H8w����-��\>���Y�#��0��m���?1��������xҀ�6H��E,D�K�$��.�Ю(�/��[����/J5s��=5 �}x���+Q�郙�ZjeM���;�.|x�fLt���%'z��Tq��^zû���hm ��ꨲ��҆��>�zO)�>�-�(���!�����ƙ�<�w�˳>���'$#}ׂO�|��J^Sẛ���8�;�JYA�Sq�&� �N�8�|$M%�<�[?23E�h-G�O��=\�T]1�ݹ0�Q�-C7�
Nt���&��<>:��N�P�E=�{&�ړm1����끎� &H���f�-�cK��^Z�)41}�E�L�G��n�q[I)+�6�(Fڼ~ָ��2����c�f�,�fS���#Y�'/��h��8��8]��$�� ����q���B��ż�ÁÜ8|ĪT�Zv��C-�{����_> �Q˓/H�����<M�s�x&�C�N���m^����������ۣ��G`�m#Ϧ�h�:4F���B����> Ú����$�����ٲ7���z3��q'\���JSI1d�����d&�#r���O���&���SV�P�d���Ǩ�z����P~��;�8��zS�6|Uy�J���
�����и3�*�o���@�ذ}!ɼ ��*��獋<f=���0�|%�@�������_�H��39�@�\�3ǣ�s���O������"�7&Z�Hk�V'^`�M+ mO`
w)�HE�W
	��=T�.�3�����l�J���)e�>�d��$�F�a�VR���>��~q��!C]��~��~��I���n�Ø�N�˷��8��gh�6�y��Ǹ�,}�f���w��Rۗf-�t�-I8Gi�o#>�S�6�������8��+�������f1q��#>4"����>���|��"$��(}O ��}� ����zߠ������߼��)�]G7�`%�����-t'��m���y\�#�B&H�L!��%��y���H!����:��ּ���A�m���80o=�P<����v��h��zı�rK_q�o�׬�R�?�E�${��'�� �7�\���<�e�?㟵\1����?��ҋKP�a([�;��9�-N�*��^��W�p�b��?�ql��q�����9H����*�����+1����lz��'�6�NH��F�=�y�8�x��;�e��F�'ᒡܨ��r,#R��NI�t�N��4x��`�\����k�&��IC�M���fNV-��m5��������i�/����c�՚�6�E���h�4o����i�1i�yw����F��-���)�6b��)2X�0�����7����Z;�������]�jn��A��T���KF��o7&����@"�h2�K�v���%u:ͫR���K<X���8�x.��|7����K�l|$G�X�"$��P�\�����n��W����1���kR�%���^�tR6�k����R���@p�E�K�c�a5�}�_o�V�Q�~Wrz����*���>Q!1��u.?�N���U8��4(;É�x���ף徥�;�0,�غ�kF!����i����%@��ET0bp?�9=��ƴAҾ���_"��� ��y^s�$�Kտ��Nk�i�"'I��xP|e��%}�*\O�E�h�]�)�o����=y �+vI+y��	��}0/m�'E����o�|�q�?����%L����_p7#��b6=�kI݅T ��x/MžM8��<E<��m��`ݹu��P(�gw���/��Zkt�[���'��{cq�މ�5�B}N�Z�OV�L�M���ͯ�K.}�>��_�yt�<������e6D�.�F�\Q�bY�8�`����q�k�L�H�ĥ]1���E]�B�G�Ѐ���h��������3C��_@,g����#�^�#����ž��o�����c��.�CQ�裋[�� �Ö������X�&"m�"Q�;�L՞յ˿Q���q�.�w���2'��ǉ���&�H���8E�1����<}�Af./;%��v;D\0"�>���). �8���Y w���1@"�|�Z����G@	�OSu#+K7]���z�(P\Ғ�@3ѱ�!G18���!��u������5P�����+]!�'���2�U�>QZ�`q������T<D̓��Ⱥ����{[am�.Y��k(^V>O�w��_Ĩ��m�����Ϸ.�%����Pĉ���Â��:�x[6�nT��yX�S�o8�х�f:m��ێZ+�n����!ö`b��郂I���܎�NW�k]�x��b�CQ�>����A��n�C�M^陔��:���A��bDa�߹��Φ��~��
}M���6���u��l�[�/��%%=-'�;�q��ϝ�m*٦w|%*��s�S��@Ʒ���>��+�HPJ�����|)��_��w�i 6��ib'��6J�*�Z̞���ү� )����J� ,���)1�IxH' �[������j�3L�A���ݐ���ᔃ�N���פ��'��X��,/�S!|���>Mez�f�Um��� �8t4�8�X�T�����26ܱ:��9�J�-[(ݜz�N6cx 8����d� �j�qWɎ謉 ��B��e8:w��C�lut<�������Ed�j�Z*>��և�2!R�\Er_���]D[��V|B:70��>.���5�Ó.,�ۥ�����ɑ1q�+�����H��Ɏ�@8r����8��)�ii�\�-�ُ5&�+,)�L��	��p���$2j A���S���'�G[�[�i��b詟a���$m��q��8��.�f�\��hJ�����H�8���#���SVr4�����N0��<oF�3̾�TW��r_��v3�{�`��ϔ�ϛ��ǿ�&�.�7'y�/>q�އ�@� EK��K��t�XZ�+�>�Lyq�G|lR#̖H9@���p�!�C�>��j��bB �6s/��H���PϪO$����a�Q����`�D�xLe�ʧ8��&ʒ�g�͖��<�8oa�t�n#�����Kڮw���;�ME�%77;��ef�e/���Xg	{1�P�k>�5m�L��<�WeAU�,+�Ո����-mCֽ�O0�5a����6??_j�����'17��ۀ�8x�"���)>84�]|��Θ���x$����s/��'|]��bF����|��x���&-�4���<;x���z��jbN24�t��p��FP4KnQ�)d���<vs�C�Yf;d�A�v�ʷ�Y/]��GG|8��cF;�^�c=,�T9����$0u�ZJ�~:,�Jr�}|o�<S�SL��Dt�(�1�]�7�ي\鱏�=��/�7,w9R,��b��>���6�K״Y��@f�=����Y�IWF]�O+���C�=0�v�`�I�W��G�s��J+�BȅT��������>A*sjƐ��0xA��;| ����x#�C��V�C�*�ƫ)�.*%hk�'J�j�Ba�>��[z�tD�,��%�N=���&��_�-�$J:���ze��E��?{��
ƀ�+�
Uh�=IhD��`�#8����eiV���8>�[�� P֗������5�~Q�0��J�j�I#HO�f�a{�wV�0T���3o)tD�C�c��&��q[�zI��bQ��(�d<p��,������S�����GM�S`pf3�}+��>�E��Kd�/�Y1�n
VL�8T��H
�A�ߎ�GЃ�U�L�ML�M�M#ǫ�M�U+Y�s�?�L1�`5��^Mp���փ���O��6#��-�qQ#�H�R��=���TO@��ܮ��܇�tw�ba*�89V�ߒ��d߆�)�ȓ�d������B����/*��9U�ׄ��m�p�f��ޘ&̓Y��1�>��e�V����M���~(T+����	o`B+�I�07|C�{��-)o��`�c_ ������ݜ�=��@;F�?@w�ֻ�ȑ4����!�TI%�0?��h:�[��~d��ߖ��6O8��7C֣z�?z�R�C�=^��&żc���_ĭ��7�Ij^�z�Y�Б����ԓ���r��:�g��ʢ�\ㅃ3��`��ws��W���Ƚ[l8zAw�ibs	/��6��BV����c���="������$&Lz�L��z5��Ky���{,�/�ol�rw�����o�ߙ]���@+49bǶ��6�-��4�3z��m�<�66󖭧o���>	�����Q��P�ۮ�+�jS�\5Aܿ׸{�/&�3L����r�9��OӃ�t+(% �L����eFm�~r�,Q�ߤJ\�Ib岫�=.IሐYԘ���b�c�����!n�%\Wp�5}����깼L��U}�w�cR5�`�$E�:h�) ��<VL�W�i�����r���r2�����Ae��ϊ����C2V��#�%0�'ӓ4��Ҫ�z�����P��g<>«�J�Z�R���`���	�@�,�k����=f&��`d��E��"����b���m'�X1c�= ��Pϱ�ȦZA�������B6T�9�G��P-T
զD��be�D��߻��\m����5x�-�v̧8�d����k���hN'_Y*+�`���p�ϧ��0�u�*I�f*���t����/2"$�z!����sN�#��k7��K1�h�0V��������5e��E<FsSe�c�o�B*��+�l��4����<B��	Aխ��#�ݛ��fe����Ϲ����g�s
�BQ:��̰�O�@ z�!Y&�����	fܐ<����󎛭��;��@n�3�N��cJh[0��vݨ��\��tR�B��~�1֪5��ZԨ����8��A .�<�7��}��iv�������:��9�1�F���I����wؐdGQ=���R=I�1�?�Π	�����A��=���)�d8��&Ōv|�><4��Z�����ɒ3s���Pqc�ptaA$l�\j���W�8��Fr�STʵ�#�/)�Ǹt��d3����`ڜ�]hQ(c{�����z�}h�|1}v� ��(F����K��ϭ`��n����s����]�g�XL��7�5�Y��,l� ��ʙ� r<�}��P�Ci͚�E��ǚ���kd�p�wW9�Zs�:��o$��u��7/��iM�A��3�j.[��=�TOm*]��!=б������ó@�'�wXO;X��1����7�j��w$ÿ�gZ��f.'}0v��W��0q[t/Mr�m5��T�����TDI�zd��p2ߐ���\�ᱛ��<a��tU��Z��³��	֊�VV��N��䨔�"���c�����؊m]$���R|�Gh�|�W����>���Ҽ:�i�4)�;�̃ y�j�Ƣ��פ��p�VI>WH��+ `bd��
K�ŗ\nJ��������t���QI7����͇o�-�h���tU|{���Q&��Yי���<,6����4+���~�IÑuT�,��� �*4���,>dx�����M(�M�r6��#˓�1�1 .&�j�2W�-K�	c>*��&�7{HS�W��)a�����Mo��`o\?�������6���h&@��)C~���ݗZ�����M����C?���!,y Y�?=}P�D��k���9UM ��D�]�C9�=��[�Ԏ	����w�� � ��d�}Q2���ڥ�Z��𪳏4�y�s��T���<z*��-��݌uV��%]#�����qr��E��~8������/�����-SE�k����}�qY0�I�R���A>>�`��I}&�1��A��� z��o�+��ٶ���nG���;���Z6��79��cCI��#+�3G��:ދR���h��e8�`�	]�0{,�5��n̑c4���p9ϱ�v�k�He���~o���bR`D���ٌq��yt�B�\/&xϫ���I�1h�ժ�i�L�b��3?p�W֖�P�yb��މ	��z��� /[ֳ�{��� ���� �=���>�8�xD���¸�ۣ��m#�K
���-(R|wLz���yO(������5>�uw�W�=8E��Z���p�J	����TDo���\y��LU1(��=����b\��R��"88��}'�w�]C���a�~5�+�!r�Z�ĕ��IƐ��w�����H?3����`�
ӃI�>��,�Ձ�H�W�t���C���4��F��Z��x�(�W�\�8��\��g�.0�#L�7J}������k�QA��ߩ��m��a�U��������&1�����|n��9g��q���6�5ѩ_\y�3���C�B�ۥ���iab}9"�YΧ�&2��2P;{ �獉��ڦ-�d���~�)f���O�{��ז���ə��ih�sB�5��$�ܢ���7�fjn�C��(�Q�s�jX��v��WQ��Գ:Y��i���m���R��~f��JX��#2�t4���o�,6O���y���gHc*U�"̴�a�=۶cc�m�;}ӧ�<GgJu�Zm��j�TUX���76�]$I�ኪ^���,��%t��Ǖ�i������<i����qq�y��y�����EX(�־��)*?{T`T�¦�#���"e	Em��=�r1(H�G���g�VGa����%"�9�4�9=r9�#�$"d#���2���'����.�\�z�ly3k���u�m>�[Iҩ�,�Ĳ` #yݓ�ݓR�*nL*;��T�m�g��EU�TX�9(��%��B$o�����%���9&��y&!��c�Ō��~"��O�V5�Gw��}�%l���D�o" �{@�A+ߠ/��{�pY䁲2ĭJ�D�����1rY@���1�Խ7��@��|&|����oq���W�����tU��C��#���Dr72�4 RZ��q68ν웬H���F���/��!@s�����bk����8�6���}>-)(p�p->wŌ	���n�dO�W�ҏ�u`�^sDF�I�V��٨sȷ�&�k뮵]���7���H��`��܎�1H1����l�gH�6��U�$������֒'r���c�7��*]n�
�]~9~�����Fj ��_��9$Yf��
֠7"ܡ��c �
�@t��Pћ��,f���wn΄�sN<�o��v����ן���8����Wl ����h�Q,�q�n%剮"��?d�n~/i�~��*bR���jxqs��nM��D�cc{�ȸͫ��+5WH�$�85��C������1@��Rj��SXo�8���=\�4��a�^a�b��@I�� 0U�_��-��֭��F�3������qL,M�F��V��w�s�<[�-ZI���\N��!S�Z�}{�����(� ��@wX��Yx�?ˁw�GP�����[�p����\�O��lOzʨ�8�*�-��Xw�L�.���Θ:緁�g�~�/���>�|�̏2%RF3�5��i{ۄ0fQ�;�\�=<{Ib͜�����i أ^��O�?1�q?Ҧ�q'� L�������Z]tb̟&����F�
o�V�<���M�E��n'���KPʲ�W��!Ǝ�`���(�t�}(��)�W)#��X
'O��:��������~��>��p��y��s�rR02]l���0]v��qÝ���{�3!ꋢy��}�7p��g�%� 5�!������p�����Y<g-^�����b�� �]�9��;��x�g����-
(� ~�}�yS����6�J�#�Q�����K[�z6�va���2�:A �7gF���8`e߶܃(ͬ(2������hd��He�JHHSJ:jU~"щ*�"U�m�̔�!S1��#� �c��C�����%�������q��زY/��*���Y���R��T�X�s�|�E�1fj�u���r��2�������=��o��U�1� �ʣ ������ )^����[���!�!�>���}�k\.ALZ�(G���fӡ3��u&P�z'���hq�	�s� ����S��|��n������&�&� 7�{�EK<7N��F{���b���ԳRL��D���t��R���ٜ�w�mvy�@������Zu� C&�ϥ��r�3SAn�d�S�Oǀ:V��'O�kƉZ���joEV�F� P�̖W*&���؆�|�ט�7Z�<�Ӑ���J��)�������+nW��7�
�t�������j��aP�R�z��sh2x�e�S���@�/��jB�q�<��7}���}���~M�����G�ܚ�X�u�;H:*�{nW�����~yԝ���iǉ���p:|5g�����}#�� �E�o:�o[�C����v�ה�S��������N�꣚��q߉�O�W��,7dP��߳F9��	�Z�q��B��a
A�Xkx��]�}07�㪯5"���ZG����Qe�fG����uݥ�=-��GdhMF�"�$��ԣP�/Х�L,��[�Ɗ7��d�>h齥j�;ŉ~�dK7�B�Y�wu]g���B����ս�ŞV��7�Pq���
��\%j�u��6�;��htWy���*^U�G,6R��時ŵNMյ�̌��WF�gʢ�J�?x�1G���RR&����gZ�����s����uj�WSU�b�c��D�c��DG3X.{]�����sM��}�
7��Jy�3�|�F�X�^������s\z�x=�\g`�8S�Xi�V��d2ʟ��N�	�5;eIr;e���b�Q2�R^6�!�����o�+R��t��Q��R����\��p��:K���C���h �md�a2��[l����Z������s����w�㵪���	TK���k4�c�a�@E�DYch�> �\�e�L���szp�V��Z�ׇ�\rÃ���5��_ �`a64q�T8N[�sa�tq>v���L����8s�R*��O�oޟ8R���ptԪ�^" �ڽ�"�*.��ۊ�<�$�
.Kb�ժ3�
%�6����t�q����!:�/=�Y.��99^<��ޛ|>��H�� V��9m�Jnp����o�7����Necς-���Lh0jz^�5�ָ��9�6�.�a҅����á��U�i�Y�5/d��*�}n�KJ2Y�Yԋ�/,D���t�G7*ŏ�O/����z�7f�Μ�A��PL)��,����S`R$`�h�q�qK����羚 �*)=C�/2 e�Yl���yۄ���bj4��j�'Nq�̏���*���t�S���j|%�v��Nf#��]o��IH�(1�Fdb�5(��[�~�ئ�h|Lpx�X,#Ks`�H�<�X��&OHx�ϭL]�g5WmX-W�͡��F4"-���6}~�̝�Q~�F�Q��U��ݗ[����U#�׫a�q��ME��GY���۬�����H��M��E�Čw$�^�V[ԗs�.��И��m���Z�	���׷����M�l/G
w��!���,���"�Vo� c`�)d �"�e�hK�s�V��׬7vU�!�_�w�N��Ry���[1+�k�>G�ab�z�g�P��.
���3ː�H&�j�E�&���f�#�enDـٌ ����{p��ؤn������/0��o�������tT��.G�&o�U䯰�w�n�19sP�'� 4ڙ;�T���B"�Vq1�#�P �����89�F�ZΧ߸Ԉ��	�U4�� t�߿��RKn.�-�����$"�3��&��I�(�9%ə�;7�Qf��4���;ϙo9��D��@v���s�፮�\�$^T.M�g$���8VO]����K�J��"��[}ws&5�Ɲ,�o��;���r��qi��"0us~�h���:�=b��w/�����V�!�V�����,�S�| vE"�^��J�y�H{K0�L�Gxï����>$O�=�3��?ػW�vvVw+}���G��FaM���*�)���y�_�����\I�8�*��u��KF�%���;�9�w0h�p��gpՖo�~XY��V�e9<�m��V��ߴ�RK����]�z�j��jj�+/.E���CcuU{���"D�<�Bj�����"2VTczp�]E����|�̯��S�[=�m���U����9gwv�(�3{'���X��PTyh7��m~Ԕ0s�-��*�_ə�g�EF��� ZB2I�R|#�����gI4�=z4�s����҄�;�}L~t����Z�H�1��'lo��@"'떻�)��/e�A���=�d�(b�.�/�(Gιt?�=�[�(Ճ��`1AT�x@���bz4xB��U��]�X]��"Y<���o���� >�FI�[\t�IǤ�O��^�W���G>0��=T(����ω�XG�!(^�@��;3�I޶-Q������@��櫯o�5�>e���beE�r����<*��e#�8[��H/� D�J��*tKet`9%�9�j��a��|�M�DpL�D�F�Iå��&�s�bB�B�ₑ
HH�iR�&��|���f-���?gCL(f�!h^�8�GY��ú��)Ŭ=��G��;l:5ղ�.�g.��g&yG�K6TQ}FFԙ�d~�����h-����'��ͫ���3������2��3����^���R,�SE����N4�^�8�1��b�	�����4������ yup�!%�>�{����ŧ�7�t��uB>Ξ'1����<�Hl���>/�]�N<���/Ͽ���ںX�F}ymR�澓_ۢ��|f��y(G�E��;\��ͣU��VH3Mb�`�y�����x��aa�����X�Z���35�}�DRLGQ_�'F����?=�ҔMo%f�u�{������q2Le�>��y���N�8�pw���8$[�y��>���"Bl�u�0��v����R)�����m>QԬ�hp�랓ڢ��O-�gϞ��"у��%�������R��K�j���X�F�*���4,��)4qwb�X�,O��v{7�UVo��of�U$�>�5x�I�_L
4��>{?�=xi�K;�f#��Y�htKJ8I.r���=����]+M�3osP����ƫ�5�Ùq��Уr�i�^IɐK�f�w��EP��$����:���2�����Q�aY�$�G���%d X9�>+Փ4u��¬�v:�j��l�P��S���?ݏ}��.�X(~��Д�8�Ϋs��W������Z���VR7��&�q���<�,k)�W��j�)����~�r]33�a#��4��n#;;�R%1�R�c�A�H6�m���󊊢�w����vT�"�f��^��>����2�ޤ*Qg��>%�n��h�v�����t�P>G�z��WW�B;�k"�
����ecsSV^~�`����|ck󏵫�1 ��h�Z(Gn͈��ͫ:w�w*y�y\��F2�i.FД�6�6�{��/%�/+�kyh�-_����W2�+�����)�=�����I�ڔ@��gC�IR�:l��0��1��1��^�r��������B-z��A���ɉ���а��8i@���D~n������G-�}>�������g���uA@���gnll���,�U���������8�C�w�ݴc��PL�	DO�8
�Uϒ��5N^G�q;��t}td-�q��CU�@[͢q�ҟo� Τ�Q#����c�|\���5�{�����e����ܣٳ� 9U��GW�m�N$,�����M��5��-A�=|0�2�L�-��- @��Ծ�_Y)��bܠQ̛�x�ug CN[u4�S��4b�^��c��F��>y���+�p��e��Q,��1�jĚ�Xm����}�=O�]8Oda¯�w��C=�_���S��66�4X��F��;*f�oq���E{9�~>�;��{����o�m~*u�C�t(��0W��ѽ.��w%��2��p=��u���<�֌V�񋋏���L�ԨQYQat�گRgπu��5NU�ǣ�&x䥥�rrr����.�P�Zf귯��I�rǲ���I V�I<1QKC,x�Fv���O�L���x��^��U.���)-���u�e��a�&�,� M�{�3���zyy���U ��w�wf뙹��8�':�5 d�2\����Z�U��_K 2����7V�^��肬���L�͵����r�bV���*?N�b<� _�B8�Љ	CLǱ~��=����"�(Tߖn�	P�?0L'aG��R��Hzt�������yu���9"���%�����ѐ:BO�b>]E��'V�ܻ2�����̦�� �&+=�*��l�j��U����+KttY[g_ ����Ll��j�j]��e3�V\u�E	�+�9,]�U��h�Uc�fp�Xa�χ�)�HE���+����,�T�����G��s��u��\�e�R�*ʽa�q�E��gnM��Ԣ��/cm����s*M'���~���Ð��R��(�B����X�.NL���z�h�aο먊'򇇥�%7�Κ�Q@^0�j.=�}r��o(WK�X���*��1	h�a��-�ᙩ�Ԗ��(��F ���"+M!���*��dޜ3%u�}��ȚՔ����ؚ��(��.S�fʶ�$�������Яtܝ����4�{cۭ!���o�/}�� �2l��j�΍s�>�v�����H���93��L�X�P�,��,���Q�E�Z�f8���И�ʀ����K������-��2�����/�H���L/@�n���U�|*���r}Z����E�'��������w3�����I��΋���ݕ���#d5d x�S�{��1���I�H�k����^=�1��hCM��7�(R' ���SS_oOU�mE����zz6��&�WY�;�Z�LsOy;N��r1���-�QSɌ9�'���������!�-�\�('gt�1&�+& @yzz:�N��Q��!�
�D��Ӓ�My{�ʼ���37�Z5��5��:�㉸g����\�t� �$g"��}�T�K���r���fE� T�7'!!y�]�j���w�����J�A6q~��)�`���??�8haw��G��@8���ժ����|��`�!�����8�>�E��"��^��p|��xb,(� ��Ĕ���#-T�41�x-���if�������Z?>r� ��읟���������; /���ē,^��\��\���5�������Z�/Y�W��>X�)sG���������J0J����r��O&����t?��JJp#Ї�	˒�|/ܩ��D��L�>u��D�0��8V�d4�����j����.�R"�+gh���A�ѠD���p0��R��@�>�y\򅌼��`�f�'ǜ)&�ou��o`>�7h�m���gk���� [\�sx�E�+��y�<!oU?�H���/1�B��LB����A����Ҡ
F
�
���[)t�4����V�"##��t�� �212�E��$�)hjοx[	d���[".���{�
(wu����9�ɜ<�p�����5`�w6-�����'B�x���*����\���܅���4 ��}���N�c�	 �� �/�f��((8Ck�n���ϝ����l�O~A�)bA��]K{9���N�\�/����K��Cӆ�_�Z�򾮝ݡ<����]���D��z�~E9u�����rTD!�b�L���z�񩕬zƶuuu�H��c��1qqy��b�~z�Gc�DKǒu��Z%�?��6�(�����ʛ~�,F>3~�eA� <;����.�q���r�T'p*k�s� ��b��ū���^�xΕvE��	����t��j��lYYMM����a
�4YGG���(#��R�چ^�0E@�}h����;t`u2�YY#~�L����>���3��wp̶�: � hߙ�V�,l�������0	�=l��b�E2�XXȅ�Ů�ha�;H@E�zG�b�W=P�`���nM�撈F~p�UH���);�4����-��,�;t�9���m_ e��]3r��6���4�v;F���dPS$�zv�L!���0�F'_u��W��B�^=�Rk���C;�'�b�Xܵ��,k�d�"�y�Ga@b��m�i�y��b���v��(y����/����.��C ��AY�::���7�2Ĝ+�uV}ӑ<������ �T؏q��8b��%bYZ;��'�HF0 Fʖ��dՀ6f�K$.A4l���5{�BۊWp�VV��\��\�g�SV�pl�.&�3��Y0��2j<���@hA���;q6�~ɭ�<j�F�S>p�8С3Q�g�pfE ]�d��+C�.����Y�����w<+�^d{X�?�˴Ҁ��� ��&R�>�'�������ʵ���2��w!N�P�ra���N&M6&�Db�R���L�(��4*Na�j��	��x�o]8T�j�aa�)� �]��d/`�5�.e1�^3b���oQ����7�!�,��F3�{0��7}_��w�o6Ζ*����[�祏�#�"X�c �b�>��|\Ck�<�	��62��YI�,5���]��Xv�V�҇�n��Ÿ3�+����PD��LvKŮ��V[<�J��l�y�������M�r`����F�j��+/5��k��d�y ��|�򾛹�"F��v�ɴ?b��X<_�}��Ӭ}�	^���BH�}�G����bP��|R�K�a�֕�_����)��e1��:H��D��@`P7T�����_(��r�[o�2��H�z�%�ti�񼾊��������y�Y$ ��䚪�Q��&[����s��ރӺ���>�����"���EM�NI�����b´���!�v�i���:�ʣ 3�A��P��A��Ҭ�Q�淁��.��,���鰱��i..U/��K�O��h��v@��4��^«�i��`9�Vm-�d��[�S76d�d��˸d$u�Id�Ӗ�R���'[��1�f���/11��қJd
A�8����~��;j��Z:Ȱ���b��P_'�{[<�t}�1��$�m�(��nX���4^��N����M$�(� FM�=��u������8)��<�k����mSذ�|�3&Xz��ؕO��ǝ���7��〳��EH"�l��������A&;����t��[������yO�Ec��x��.�	D��QD�$&�#m��ӗ��Z�z�	����R�q���]���C�$�߹͗s⤌@M�����Y�quF��"�ݨ�@�~ߦZu�Fp��/���� �g�6�b�T��J*���i��ً�1������O�<��C�����*�٨��<rN�AkY�Ga���a��t&Ҭn�=2_E�;�����0��V$��ؕ���7x��� Y)����\�dCڀ݃���ȷg;| EY!��Ϲ� 8Ņ�Z����H��	�����ch�jY�d\!������zX��7/DU
��?]d�`��X{����%p�-����:�m�i��	8$ 8y��f��ƴ���E��?H�� �!/޽�e�G���I�^l����[oJaE �0�K���W�o��F �P�?�z8H���\n� il`l������Ұ��~`��my5�C����hƒ��6c�����J��tv��),~��̳4
o3^US7��[.	Ս��[��������Cw�X]�b䙩B�����T�Ze����?�im�J�V����<k'2wCC�(�=$��!"��p�{c�8�v���D�����D���9��I�WŐ�t�������{�EGQPDEz@E�NEB��A	���PBʠS�F�C�Q$�s���9�E�~�ι�u���?��wV>�y����Z��Y ��e���p<�����кGyXoB���~��l�K���[Z�.�l���36h�!�?t���%�Y����b����F{M������|Vx""�daj�Ra�����(&����%�Ba0!�m�ۻ���"e��+�N�(f*��L(������E��G�+������/�G	i�?�qtZ�+��y�#W�
i�rTǍ� 4���n�Xlۑ�������x;��EInc�T�뚮����G-�a��9�j��F?p�u/B��*c�!4t��Zy�#q��ġ�G�uE�nFY�2|�u����ܭ�n����)�J�N�J�h�������_�}I��.bH�yI3mM�b�a ��ґO�R��$"ᅫ-��~�쯏���>�D��Y�|s�ʧ����c�h-B{e��AFI��y����Wo�<��T`��a^�M��M��)� ���U��4'�4+i�گ{bu�f��-�Q�\I�m�J�<�g��a镴ݘ��b��[M�8����݉5ǗQ���!���7+��h�E'(���S�5{$�	Q//��p���t
=��\:M�|�Z�Au5[q�ar	�=Ɠ�����l��"��H@��<U~G�t�-N���"�C5f�r�?�f��+/1+]ݫShx�-~���7k{v�B�<G�wg�-v���:���u����K��%Ɖ���U���'
?��A��s��Y���b���ڪ���s�f3��jL<F�w|��V�c��B���w�'�yO�����%Jmk�a��*���We�#0�T�!�ЃS�0��)%��[�*���ڵ�$i�<�G�Cr93R�r�Mp�a�^��>�oJE9�Ђ�d0l�f(�����h�K�fG�!$֣T�"Oך�����n3�Z�	b�c�'��a	�x�4!�����v�vqФkȧ<Z�׺%��5h�eA7���Z~�m]V�{�◺�����>�^'	�YW�>�Tf[wڂ�j:�N=�Z�+Xx�q�A�n˱��,2~L���,}���?�O)鵯F�B�tz��$�����n[���n\K���O�p����	�^�}����!G��r6��,菃�����3����i��r˱���#s��N��q~�Umxv$���^�%K��o��.mX�Jhg�a�mckV�q��)�e��HZ�iԐh6qR����܋l]�4�m�0VO����Qe��$�Z='�M0���{� �'(�L�|��j�c�Ͷ����aORl���>=�*']���C��EZ���h��(�eh*p�yp��Fޑp��twr�b�2Ϸe#��Tmb�4�X=�����dJ��e�,���Dd����QJ�+��#�ۿ�+�5��^;�7�y|IŠJr�/	����uꆗ^�'�P"U]g��ֱ����$��h��L�`_��I@ĩ�h�K��1#��ۧ�2�G?��hߣ7��0��m�)=S�5��t�'例̓��1Q���CV5�Ѽ��z&�������[�5���ڄ�f��h���g���R��\�
�?���R<�]�����~�/3=�W��3ꇉ�
-�-Y�����Z��J�G��1m�>\Ee}��Ax60�w5��_Z�ݩ���J��;n��@�ײ���x�"5�9:�yBB�U��)c��Qܚ�L�y�׸˸�At�b��TR�Of��N��W���NDx�<�SJ̭�Y���"<���ݤp'}�%5Q��)�e�OW�y�c�jz/u8�c#�����[��_�kH��x�[����J����=8v���å��Ƹ-��ʾ��qY�PF���c�\* ����pO9q���_��^��or����u�Z�B�{���$4�G�¼B�@�q���Q���>	���.��3`�_���^Q�?�&"��>Md����;�,#x�|��,ʟ�*��NyZ�%�r�g9؀�b�aD��Q���y�bQЂh�C�~Nֳl�%��v�W�!V��wЭ
��` �#K(G�}�ȵy������G�@+`XAG���vka�_f1E||��%��t>���]��ފ6k&1��v�����b";���+G�5ic�$��)Q��yY��T�V��M��) � �jJ O_<�Y#0Я�m9����boc��~���_���p��y1�#�S�Ƚ�N�t�5�*�n�3:\�f6z�d-��U�v9�z.Dx�;*VS`ף���^H(�俘�D�*���<.-�&6�d�#7�o{���<-�<����N��M*YS���`�*�
royA�f���AU���ه���4�+�0�G��~�Z�$��������.Y~�#ߜ"N���A��qm���mog��i��Y�3H��E�`B���/uA�oo�>s.4 :�e����.����Vrԛ��-Xva��l��Ջ����K�W�7J�]4��*���N���v�`Q�KK�q���sU8Z�U�_m���k/���4�!�1Kk�Ww��,�	����N���`�cjo�i�Dy�ll���m>O� �_ �tG����~!.	��^:U���8���"d�wўu�ǋ�TؤIHRS'1��u�� ���3��,��i$���<ܶ�Ͼ�[)N]��*H[v#o��_q�ș1u����:\�h�vS�Vg�2��ݩ��XZQ��Mu[E�%M���{�~���o~�KH�!�ӵ���
��O�ݨu㬑Km�L���_hA����{�h��i�˖�ss����po�g��;��C������q�eI��V��ۉO��|'���C
+Zn7́\(|I%�jB���1	ƛj��^gSD�n)5��DMI,G���Y��9��,�ʍݛ����I��JKeB_��R��+�nÊ�[/|��d��o{GP��9ّ�ٽbC/���c�7� ��('sR'�������B��"�~���g�槮]����l�q����ڽt�ldp�u�[&Y�Aݾ�x����TԐ�j�Fq5[�7�����X��<��8陋b��k�n�ux��55�!��=��wh�2r7��J�l<�ҫ�b�b�ᗲ�_�޻��?H��Z&� �Z}���'�X7���dxΥ'�*Ñ��%���N�����N7�9*f�+�������m�������V��&շ�7ܢ�A�r&��<�T�a�w�!����s{>�1.��0
Yci��z��cy*`�\)8�.%ʔ�t�R�í�K��W���4?���-EF�����iO3�&Ҝ�5{Q\��~[��B�;���b�cq�	.Sg�1:Rh���L(�{����5�n�T2>��\ވ-�˲WĈ	�B��0��l�N
}�K�IG{��������&��:#��� �vE��T�^�{(���%l{�gU�mv8�Ġ�9���K ����=̲j[O*O���`O�]��H�[��aNyFe^���ђh�%J1��bw��ҏa\����F��6]�U�^d�i?2P�;�6T���\~Q��A��[�`#ϴ��� ��� ���<�+��^(��A������A��e����S35�����Z�|K�������Uݔ�w	���(����5�r��IpU_�vn��ޤwjr7�}'��K��|'G�f��=�7��F��/|�k�å/쉚J���)����ܜ�%-��;R�P����|����(��0W>b�㕓��)��f��=F��)��u�2�>���^�>?�D��T����#wM��ՖT��ڃzkoS'tu�qBD\֔���#�Kx)�|���ek�9����I��Ҧ*�d���ÏFz������fT��-��{х� ?��ȯ�����Jo6��x$�S7E��+��u�����X��{���s")|"�2;��T����v��+6Z�E�"f�'���nrCw������b�K\�9i�B�S]�+�V�Gd�O;2���kZA�'u�)_��4��g�n}��D �g�I�e�0��M�1I4�p��I�eXRKޚ
DM���tm_�nS1���G�G|�3��k��k�Ρ<�Ke�z{?o'�D�H̳�g��{�P��U��fq�=\3]��q��l[�⫟9�?��-=��x&L��in�檾b�X�z�	J.۩FMrэ�E�U�C2g���(�d���͋g4�oN?���\�򾾄̇�r��.�O�ѯ��,Bf����X�� ��{h?�%%	K/���Jh�K�%C�����D�����w
��I��w���]��oKf(Yt���,q����
˝u�+�W�F�sI��2���>�+y*3Di�������'��$%~�L���F$�>}z��|�$�ǳ���uE&Z�xo2l���쾪8�	fy�"W��_�a���V�ZD����
J��w�~�NG�HcV�Y�����I^p������pv��l��6���!\�Du�O��ՒZg�e����/�DЋ5q59O�>5[}6����#Ӊ����t�dwh��eAo��K������:L��N��S�p�?E�JJށ�F?�?X�lS���!;#!���"h�a����jώd�4��\7��ao�q�6M�PC���Dd噿�{�]E��R�0,Ʋ����?��ئi�V���O����s�Tӕ�.Q+����ކ��p��|��83{��_��uY�p-{��)�c߲yt7�����^┱�6k]��J@�3�b�r���ga�"��������(�"1�'6ؔ >"��y[d����e���rG���y
گ
Y��M؟"��1
�;��:��M)�T��aVA�����b��w���v&0��ѧV�5�^����D$��:��p0�'O���w����|�t���LX~L�АKX_ZN�̢�H��A]#AS�`��f%#����ѫ�JJ��p6l:��!Ƞ\,��nl#�m���%��%���9��;j������T�Q��GWj��r��p���beEwx�0��k7T��E��#�h�i䑉z��8LT�������i���BJz�����i:�����(:�9)��'��x�ఄ(��lN�����]F�=�3�$�t�^NOO��G&'i��T���e\���P��, @8 ���6�F�����#��a��:���y�V�����J@��M���c�bv��lW�����ak�oga-��i�<썩D��=��T\�������w�̐o6"�;��Ҧ�k@�h��ja�����p��5��Y
˭���}֘�gt!tOo��L>����ƦS��bÕd�SCTS�)y�Z/Z	<�"��Ev�g`OeUUU��'~��t��$l���$��]��G���GXf�0�'`;V�!�Aퟋ9i��Ftؚ�N=ƠJ����ٴ���B q�FБvg��?�bjw�}0��f+����z-Q���	$)I�~�<O���E� �z=��,}���w�2"<<<\r?����R�!y��f�9u]p�)�9�M7�,����0�"�`u�!b�{�D����d���s���2�&�"�߽4��$}��X�� ���Sn���޶�>�%f%-m�*r�e��̠:��
3Y͆��K���Tk^Cy.K�K���PRy;iz4d�~|t ���������8|�������xUx�5��H;�O��Z�`��H$��(�h��v<�WP-�nΎ-��7"��nG19m�cV�Q����>~<�'eU/�x���̵�S3�UoV������v6��H��ө�������y�v�S�V�cnX����I����"��CL'@>��`.b�Gve���[�5f��;[���>-�������̉䱀BP�@'+�L����tI��`�[no����x�^0�ki�e�|)X�H���0������Տ��D0g�❜Ȗ��ttб�]n�f��V�� ��		]x�a5����}���&�8'R�������s��/L�r�j��bU��s*�	����d����K����03_�U,�G��h��]�����F�&���`{5�!|Lk�
��|���ŹFŘT2])^�����Ӥ�o��HW2�$���������A��/�)��jn0W8�Oh�r%�����<1izU��ZcTsr��e^Z^V��{Vt{����U��-�����_�"Շ�����[A��!�u�Q���g��yZG��Ь�ێ��$n��Dɴu��'Bf@b�+�ͻ5@���9����cώ�Ҝ��^k�.�]�a�"�=���fU���+��ɒ��ߖ-w_���Ͷ�We����q�p������d�yh[�1�ԟl���e?W>�+���m�pϜ.�Ec�������`��j��o��o5���5�A������`OZ���f۹�]�(<�ǵw%������ȣ-����x{��n�SG�`�)Q�j�C���Ͼd��[��./�O�ۦ�wd555A�j��ct�[���f��ڝ*.:�U2��ƚW�O�1�^7[&�9>6�\.u���PSN�����Vq�|"Y򌦺�q]S�oG�|;m?�~��i�r���ԾI
��t�`��1B�B`�����5�v�j�+b?��J���ڧ ��hTNȊt����r:�vʉ�xaem�Դ��3Qª��I��A���#���N�0�M���g�/n����O�y~;���˴��w���^"�`Lƫ�L0�άo8����^Im>AA��_b�=I;v�^�����������}5��)!?�z��.=;v���O�N�j]��f��7w�2ڀG̾M;|��$�q�x>��j2��0a6zcg>]�
W�[��|2/te2�u`|�:m��i��TnpHy�p�W��'y��EI�spp\�0A>�v�ʳ�cJTEn�W�O�&�}��o���h^#@���q�GoXU�[�o���D��0�������h�8c��n��r�~��Qo����S��4p%ʑ�;��5�gT�iT����L��ħ�<M���r���nv�*v��<���i*A����Xٝ�	-`$�F����$���~F���F~[C���f1:�ݙL��)�`P���g�m۰S�Y��Zk�*��F$�۹���J�-o��9f��G<�(;U��s��0��y��x�8�F�3p �Z��bۣ���U�p�!������x�m���'�Պ�Y.ou�����LB� �%�]!�}59������Rk%�1��hg:��V�0I6t����\$-�I�*X�|#�r�~'K&3'r�d���G�C���ˑF,���3��_�L���)���~���?��ڷ�D`�w��ٟ��w/��l��g��i��'�g3êZ03�t���͟m�6����n�]�zO{�W��7gv+{%��90�vj0HHq�����Lȱ0�%Ƣ�S���lqmM�\5����������J�����T�r�����yF_|���_�NA��ct���z~:��s�Ð��g>����砦�v�ch�¯�V�������9ݺa��BQ�Mߺ��Jr���y���~B k�%�ph˯�Ӄ�O������S����Lܱ��`~��c����c��6�p?�3�R����s�!<c�o�^�lw���K����1S8/��S��aT����k$'��EP	�H�R��`j�>Tɣ�}�����K4�L���كb�M��pG�bUw���$�	Z��A���5�&	�D[`!XH��c�˧{�� ��d4cv����K�ώL=�8<��i?8�T��s�zw`�w]�(kP=;\���z���d�//�%Z�!�eqP���W�-.��t����56��vm(���r�Ŗ�n
��6Z��7�(�J�ђ�PV�'��Փ�q�ޚC�Á����������F�ӃuEo�]�*YC�J��1
Һh�ç[ǻ)͆Tv���p�[��zl�T���B�o>US�r���'&10�⓽i���U���Ǹ��v�H��xA�#~]D�OZ��q�\����5�2^�ߗ�P]���9^=�hd�Z�s8�CT���$ %�qa�MǛ�7( �Gټ=���R�b�^������`�����?�9�̂�85<2Y�@+g�I1b�Ǆ z���҅�D�/C�6�����r�S5����j��W���z����� �˅�y0����m�BC�����P�<��ϯ��[���b@���h�s�E ���|��w���;��m�Q�t�Dtr���"]kP�%oP���_�Ȱjw����º���
@?��N]�S�� R1���B����^{+��M䳽*�b���O�c�{P�Z�o�T@0F��LƮyF{���t�j��-�=��o_��^ר9y�eD;��8�v�/2�y�ÓMs(Q��U��b�	w����LDL��eG8��L�F�sw��a�\	w������H,b�Z��&T>i�� �;�T��'�vui���;B�6�q3�:��/n��j!���P�B�Z�⺥�A��kz�O����!����΂��S������u��f������UWVV.�l�'�Z�k�����ېs�H쫪�x�Ֆ(�0;�X�V����C q���K��@W�Fo��Ύ���t�˯
��؉���� �Ip�
(�'z�����b�B��P��Q2��rrr�����ݼ;�,$��e @1mH����_��f��hj�@��!��=Ӫ'�������u��6 $����5'��,��C`�+���Q�rL���c�����!!5�>_�$��H��ar���M̀�2�A���Q���v�D�I'�1�C%a���tB�`��1��i�]];%s�L.a����xzA�N��b,{��K@���[.�j��Y��b�rv��'8o����A}�KO#�eWT�_����.yw��9�	Lԉ9�~��)��k�$�(!�Z�HH0O�"=��n<;>>��@�F����K0���5o|��D(;��z�,��ȣm��h~e2�C6�>�N�\����$R(_��$>h�rl���6�]<0�=�'�������U��4j���1V"�MM�4͠�Y�����P?iQQ�ˏϯ��F:5�O�W��h�����.ؼ��s�h����m�ࠜL�f��*Op���S�Y,W�0r�=�>����!IW�V����n)���8�-��A�b�(qm�D�b#�_i��O2^�,�H�C˯$�c?Î9ZX�~=�7J�X��xω��o���Iw]Q�� wz)9�Y�nI�B�U ���|DqA�7]k-Qeڜq�<V�͒�n�8e7�[�y�z�F�d�g� ���>�m�*��3�/z�=3/$Æ7]Y0rV�J�C�e� ���(d�eB[�Y�C�,�p���3\���&t$������Q�ܷ����g'[�бrkT��ϭ[U�U'�����H�"1e{u�V�h��BoUw� ����T~�S���^��=FD1��
�2�	�����?o�k-��T���xs{��.��:�cQ�����a%��Wͮ�8Ϩ�AW9L�B�YϞ���i�����������,;\Ö�x+"�-�W;��L�Vs�:�UJ��Fe�P�S���q��.��(xN�Ǹ������^�n$�g��n־�v�c����%F����,l���@Tf�چ�h��rDw���<K5���\'дUJnyX) ��k�����q�!֘Ni��,yF��)O4�z������`�ֈ3�˔NY�$�9�
 (_gaZ��zaH����cU.BOY�톹׽��i��{GP��_f��si}WN�8��$���t�5�����~R��F����n�)���z/6���ⷬ��~�IL�*L�~(j�xS��d��t>�
���K�X��iʽ�PM�8�-���sa������v�+�)�a������r�>��Sr��L�h8�m6���T+�$-ȕB�U(�$ܵN��+�1��UV���{�^��7=�񰌞�. �ûi蠟�
Y��x��͕�z4���6��X�FF�>8G��.������Y�$����mO`R}��Y�q��49��k���EDE-�:c 	A+�[<&�0^AA��@K�x�H��:ӈ�eSS�����;v��~fP�פ*5�Q�V*�tἀ��F�*跿)���f��?⹒����
\�A%kbR�%@u��x~;�.���#��+�Q�kӣ��N+c�L��)�Oo���-p��$M���t��ܨ�o.,C�F�i�i����f����v�$�W���K��2�מD�x��n\��.-�"J�δT/�"�*�)j�-�g��ν6�G������5P�)�Ct�3NΗg�sG^N��J�5��5X �^> fZ��F�z�́�c7i��N��$���b�S24�����.q�U�q��Ɨ��?84� h6�EH�<��Ӣ�ݾl����$�Y���:X)�4]�%*R���gK�n;�0 X �B�8��Z�Ga0�����O@ܸ��Ҏ5�����mYkkkw�����Գ�|`��ZuQ���� �r����F����D�v���@F��8�C�����
�����Oon6=�P����yy,��EEz���s�oMȭ���`���U?::b0بS'��� kg&� ͡@��MY㟭�t��ҋ�G)$�yUUU��h4Z�S�U@����H�cz�K�ι
o�k��"#�N�����i���k���<E ���}|�*��q4C��p���	���ܧ��\V�!� 7 �����nS�����7��=&m� ����~����\�p8����[�A0���N�xI����+;j�P��Ă�/�nf��I��$
8��� ��+{$�����^�������d_{�
+��"�~�*��$�xCh�S��C�����'tv�_څ��ѱG��/)Lr~�Y��po�r�Ȇ���\s
#����Վ�(�$�hA��X��@��ɷd�Q��p��iw6\��ѩ�<��<$�2^i7h��&!n``��t^������7H�>0xHG��I�/��Y�~�'�)͗�sn=���'�V���6�������T	!!���ؗ�J��
w�`-ס;M7���8pL�u�R�� c�Ҭ�;�������6��U�mc���-Kjk(�\s��H����ӽL�2�������h���7!y��؟.㲿��s�<>��Y*]Z^���B0	=`o�5r/����1��Y� ���bc�d�d�<�;�:f�3g��i�����n<���H�~���ݵ�����|W(�h� 5�ԃI[;;��@ D ��/���dD���`�f���}���ަ�~��Ԑ���EO�0tn��.�O���9@V�RD�g��z��� o��֣qg���O|�30!*�`ؤ�#�H?Hy@��S��r�RG��!���37>>>pI�C,�._�4>>>�@Q������~��ߪ7��c�`Χ!�R��U�b�Lͬ�ɦ���x�:H�_�z�A�F���(-D %5�K�<��;�1/���ds���Z�(8�6�4 ٢W�����h����ĝV�"�{������ĭSz��	tB���3���������YK]�[�0���3j���B@%�]�cZ��S��0����%m]��#&>`P�b��Z���,�C���8��HI�?���4��l%�����O�:��H�]I� �?��=�I$>�8#Wy����P��# n�V~jj������:��-��h�Qh%rq`��k�Cx�gg)�0_�V�j�k����4|�\�az}�(�a�G���6�k>��Z��QPP��{���>`�꺺PL`�J�G�lqlTL�`��W����
��0���������s"��GgR�����s�hW�_n�.y�*)���$�Gz�2��e�&��/Ђ$�>ߝd9U��� %n5}��D�S��-��l���
��T�&�+Ap	����e)b:h���"YSSS1\۵R��qhB�F5ܧن�V���r9�IJ<<<ɉ&��t�� �hI}��$��&����Ny�kH&+X���4�������)'I}r�vB�>�̨��?8� ,�o7ܶ�8`����.��������R�H3� ��6�x�
9�`�I�:�69I�䋡���#���mNK��gVV"���ٻ�#Tz'3���5+e_g�ЇV��(�H a�dG��6#��� �܊ y$�H��W@:[�;��%����c(B���.-�\�9F�218Hg��e�Z��W�é��t��` ��i��B}��ƍ�͇{��O�Ľ1U�aй����QyBu�1\�,�N�Q�H����;�đ���D^����P��2�.	�],d�'m����)�m�H�fno�ߗ����I�dN�I�'�i��j�)���s�턋�hWW�m�w,��I�5���JZ=˝���D3��V�BVV��%��|K���ܙX��1�T�������&<fP��m` ��ی�q.i"w{RRRe�w��\f������v/{��y{��{��F]���^��.���=9^��ۙ=#�QV�.��'��R�^��Z��<�$�>E�=*1����'���!��e����-;�{���Ȏ"�㋄:6z5R���q�j8Y#��\�<�W���`���~�e�ƫ��/��U3�M�0N*A6T��$�&!/�B��jN`Y)��"���=e8�I��=�r�}9c���/����\�r�\>W�.r�D�Jz���}	Q�uή(�^��,��uM���z��y���^ÿ����������^��u��g.��}Í6��26�d�/���݀��s��Vi(��)-ȑ����#�HP"��v�Ɨ�{��~��������4��>�8Dv�Bٜ���n4�����"�w��"
a��p�ฤʯ蛿���TS��eN!F��_���-������sGh��y��j�����Jv��é������5C��%�5%����
��,���>�U�բ�j�՜o���<�[M�#�籂o�J[?���9"�~�+�E���`�ZN�,�ck{]�Rd�o��I���^�oWD�]2�qs�L�����χ�AS�o[7<����<�$�������������_���-T���`������VK��V��w�."�	�����a�8J9x��������|oOΔ���!����I�����8��l�x�ȅ���2{G�w�*�W��AF׃$�P$$�f�Oma��ψ_��*����Ս|=ۙ6y2۠^�?=1@�Nnb�=�QC�������+�X[v�_�.h4�K#.��rA���$][��%x`v��w[���ʅR�O���d�5��Ei+x��D7��&��4?8=-#n��'g��2�n��V�O)���5�0�2+���I�a;��`�ne*�̍ �ٱ���{��/�y�~���ﻳHm�zĐ[�n�YŐ��<O_��{���*����{o�j�Zh"l��J�QD;_7G!e|��
q��u&ǗUdw���z.jP��+D�0���Y��5!�ō}��`Y%���	�F%x���}9qL�:��XD�H���/}�߬�|�|�3�@���w�Ǵ�������Y�i�;'�h�m���&�����9����Jk�~B#U!!�F��s�!���2���sц��y�u]h����W�zVWJz*�S��&o֭dj�'��jZ{
m�9�#N��c�m���k/=�B��i���oЄ$UvO�T����L�Y�h=�Uf�z��Va��������5�l/-�̍+���3>�����pL	h�[J�m�k?�z~���F���������IBQa����in����&;�j�o�E��#z����6����;�y�6NHm���1XH�Q��-͐l/��Q��qF��	z�.�"�->߲5P��`��s#ЯR�<�VeDu�F���A���Xm}|���*�yq�9����;E�,;����h	��[3��a��G_��D���:S"�a�T�ӌoV%��������W_�	a5b��� C�R�<"��|O4�*�r�RUi����1�yؤԟ�.���4_��Am�72���|3��8�q�:��G+'�t�f:Nx�
L�$q讦�{�I�p�|�Y����������ǶG����뎑��}0{l�P�=���i����mIZl���>�:�)(C���~��t���X�:|:�Ս���<Z:��$;�7T�]��)�W^=��y���멏�����&��}"^��)'f%Z�C���Z��!2�,L�"��|"��7Z��Pu���+�/�h��d����\�`?x�,6�#����+KkW��JG4Y�ZsL�1t^?9QТ��ʪ,��1����r����~۞��S�T0|r~��������)�q�9����h�7�El��[տ}��*yd�{W��������[��gf��_|IT����L�7�^ԷY��&�y1���D ae׳��w��c�h��B���>�����Lk�� F����k�?WR�@� �ȿ�C�j�,S�r��6H�?����/�8H�|���|_�>�c��x`����oU�;��H��g�K�E�qXX;���e�(��j���.���I�o�g~�L�QI�˖�����������Ӳ�������b�F1�Y�&Е�j�o�W��K�+��mzR:t~߽
8��!~Gs9��H��/ �h�j��}.?;|�wV�����9Wo�]����B�����p
�|^����N������&7[���~6�8�oS�KeBש� j⠡��� �����]0#ݼ�Tr�DV��L����7W�`}uA�܇_7�b���+}��[�wZ-�*a�l��#͠�����%��I �f�G�s�]��zpy���|���_���/~8�'W�tf@�\������s��ۗO���I|-��������&`X�_k�i�A���F�������p� ��Qã�.
//�ƍ�ɼ�MϾ��}y<A=�!�M�d
x�OvN�Z`�2>�Fti8 �fk���.��K"�G�+�9O���+��kt6�THV�oy ��αC��7Ps��UP~�3�_^A�yJs ��d{կFD@��LDQL:`��|>�����mǮ'��V�&s&Ʀ/�^�oB&K=��{n�)T9gV����om�Qa�SJ��3��q��	��B��L���d-��y�KhW	�r�V0!�2�{YG#ǹ�r?���x>}"��F�u,�W
�[x�}���bx>�դ��N��Խ�W@{��/=l k�"~"�<�.����p��֎6?�����9�n&��U6z�C�u��y�#!��F�@7�E��SZ��Q�xo�a�wѸvz���e��ɑ�������+JqQ�k���&l2�t!?����F��C�1����!��у��(A;\��4��N�f�7��4ҰzH]u�Q��R����fa�N�{�2O�֝,�cѻ��i����6OI!R�}��}�#���$JܚA�T	U��f��^�C�z,=���2�h ��%�g�_���M�����i��e��r�b�9�I�(����C������#���~��S�G�CN��� ߔ���"2R#(0h����c��c�j�6�oͫ�_��F���r&�9�"��^"GS�XyKP�/��2�����+���R�j�j���&O��<m'��=�����&7�(T��X���}GM���S��M��GB���Q%1ڂ�_��$�sS^��Y���ç��s╶�ͭ.�߼}]��Z���M���,P�k��|�]Qi�5d>u��=��d���/Er~��Hɋ�E�/EDM�ѭ����{ ��_�8M�=��|0֎WY�|��.�[�o�c+�kv���3u[+ӄ��ֺ=J�o�  �,x����+�x!�_N  D�ܸ�������_f~���E��q�<~�ͩ�>�{���W����w������M7R�<��~0�]��:�6]p���&e"!�޵c��Ƽ��SV�K������������A'i�D�]�C�+LD��y��k�Gv��Ea-�&M���J/��K
Zҥ
s,�d��״a� E��t�n��I����ЎiX�>��D]_;0y��a2���x��;���帾̝� �/���t���09���aϓ�l7z�����G�#]'V_9ۃ�h���K~}�P�u6wGM��#��r��/��I�q�����^���*t1��k�Nz)Wh��3���-�=a7'��$������Պ�c(1�O�_!�&YK��u��_Uؽ���ba]~j
�n�k��R��������Fma��j%}����l�о�g)��M����O����d�~�U��&���c{G
����n����g��+��Y�Fv+�K�8ٸm��\���8���P5��B+c�g����RF��1�b&�0�2LH��<>mT���_�16j��W�/O���U>���� �Ϳ5���#��7�ޓ��.�e�,i�?UNm~��%�៭�4F�{
�I"�GƙP��tRfu�{�;n;X%6?�U�Y�}䇽����Ml��{��H/���B_�e e�MF�-WBS�f��<�a�9��Y��|@����uP���Q�ɽry��@?�*�0�q�C:���j謒'Hl!!q������x�f�i�dF�x��&��"�-m|��A�<$�M�����X�y��/�lP����ԧ6U=ϥp��`��C"/3!����*92��V�Q	��E���|�}Z)HԌ�sg[/�:M����%M�k���'2�O��zqXo�`�y��wd�/f�7{��N:�.5���f/K{+I�H4 �E����>�M�x��(W*q|s�y5s�"�8�p���W�?���Y�򭽮g���-�"ƪn���Q�6�.���&�o�Q_�.���B��X_ꔇ��@�)���y���Q�L�����/K[�ߢ?��#��Jk��5������	���.�D�'���#3d'�����urxsޙ�C.P 2C��2&^��Щ��+�`͚�ںC~��8r��t.Xb}9&��mv;�c�ez��)��GZ���\v;X�r�n�^��0���2��5���?Ҿ,x������X�PO��Gg��n� ����rQmck]wi̶�`j�a�����v�ԝI�"���=7.��~7�*zX�f:թ~d䫔�Q���J߯�,Ƀ��ס�{#���e��)b��!���}�Sp�͎�Br8���L/m�C���믪
Crn[�;φ�ƞ�}6Z���Aq�i ��;QFSgD��w>��Y�[ʰZ*��cUy�U����~�l�T�?�Tџ�Wc�Eܤt�'M�_R��-T�WzW=���@la����R(6��MV�l��V4Z��_V���p�J�5ub�{�Y'��5�o��\/6���M�cr�/|�I<��ۆ�.�T��K�~"�e��s��\�J��]���?h{Ϩ��vm4>��<6PZT�*�&��4鄈�R"�������H� ����(���B�[q���}�8�c�V�+k�{��.�5K�n��ЪU��T�Ի��"���#��e[$�s�wTڃ2���:�#��}�PB&b�e�·�4�4��G���J��3�)�;ќ �pP�9#�]W���;0V�
�LU�&9�bjE&�P�bS��~t&S�{W�S�w�O�{ ����z�%H�擹t��a�Ѭ�_�u�Hr�z��)���mmM���'6�1���8�^�N�*�u�^�#�<���������%��� Oya�6��L�2�zxU����cэCR�@S��B��"	�E���:^!����1B8xӴ�(�M&0WCGS���:��0> J����"Ϻ���i�&~>npics��9�}D��S���_~>*��8���"�;P5D�d�		�����B5�_C&ܣ>����%#n,j�˯�!��U���6�7C53�,���,}�ݫ��h��q���ٳ�@�+L�'ٮ��γ$w�ӌp�A1��=/<\�d��Y筠BR؊]e=�����:�_UQJΰvZ�cV(z2y))��I[̕��V5���M�Q�`ƶᕪBNb����~6i�gZ��2{r/>4�˫���DJI��sHm�C���~MB���. �0�*��֨�Zxqb
�������~]��XkщGZo�;%��*�|t��Bek�k���<$q�.��:�F�8��*�5+yM��"q�DB���HD�!��F������w�9�@��mR8lLc�:�x+��E��(*�2i�P+�i����J[^�0�\�/�bz[��tdR'�g�`A��MW�9wS��6�����U��Eb��<8�D��I��xWY� �z^_/�QaֲS����H�~�
���*��)pG�5Kǩ�4[���V	��br3!��'��i�J<�q�9�7K�7�L�X��ϰnn�'l��ډ�^j����z�Z��5��ǭrW�L���՛�%=��s�i�z��[z5��=A�<�Q�[�����r�Q��/?�T\��)�i���pI��S*,�qB�� ��}�G^ �`Y��9#�"}"��29G��Ѹ�����8���+�g�9L��H9��'�Pu;O��p��Z_��DIëFg4hd��Dm���u����l)�K���q�p0��7(#�����#� x�0���[���n~3't��+h�}%����~�18��]Eu��ID�q�鑫])�@����2��t�C�B�O���ac�^����9��G���~P�ǡ2@���B���Ƃo��]!A���΋��N�����n�E����x�")5�Xm�yCv$��Aȥb���ۏ�����������`�,�ck�(�2�J��T+�t�\e���w@1���2�u�R+{b�Dۮm����zxd<?�%7�v"vn,I�v�Jn4�z�)/y�H�m���,�E���#
��^S��G��k\�,�� R�5�9󌤼+e������S�\���Bx�3T�|C���G�(���kSգ�KcC�:��(����o��^UH `n�s�/����O䷲����B����m���Ar=�)�������ɤN�	�(#�Y�#c�n:��P�y�@���Q�������}�̈́qS��A暃Yn�'�� ��2�җIˊD��j{�9n
_��P^��jb�e"�R���KL�y���K��R�MK�Z�nB��i�D�7G��逫U�66?f	fn/�BP� :@8���������@�.�E���#��5�8�|Jf@��d��?����i>Nu�%r�����U#��6��'ɻ��'���3�F2��Z1�&1 Fov1��s���L; �'U=�[@>˽���n�>�j��%`��:�rW�r���-�e��c����n��D�t;&��g#VSҁ4�2�7Z)*�?��l�0�26���C�]_ڹ/1<�,pP��"�:Uq���i>gh����o:ߖ�����IM��s��y]eh��)��4ax�v2ǳ��is�X�S��r�*�m7RC�6�JD����N�NT����n�<���	�y�(��'�BCj0��av�m�|��?��ߋ<��uY��M~������_�d{��g٨L�^���V
�O��_7�k��463m	ݣ9������3�����l\Ό��/�����#!�׍W�!���2@���,��[Y�uoF>��x��ϐh�º���j�+��+�]���BGQ_���A�~Z�OJ6_�r�g ��� �dçßBZ����Ms�@\K/s��/��"�1Q)�t��_��V��N��\wC�%/|��`��:'�ß N��K�L�M�z
F;
8�M���ߪ{+�PU������h�߅E8WmL�����Qnc#�a�i�ΗW㎰��|5.��}'A�Q����i��K���Dr�U�L�t[�;�ڃV�ej�V��K�ڽ���CAF�C;�)��%2��^.%�v�)��Ogܾ,�.�	@T:.F4���PЮk�n�}�ܱ��������)A��ř�_��,�,��{�?�d��D0v��乔Q7���6C��x����A�r��ි��2�d$�Zc0̈��j��P+:g���+}������ϳ����k6! O��q��8�ԛ�9+�g�4�W�ϛ���u������
8V�>i#qiH\tBs��qR�"J�r����;w��j�{����p@M��s=:��m!zs��T����J0���0�\~�ɞ��n�����0z(��^� �"4��E�:���ƶ\����V�to7ʸ��4U"���g��@�����R�c�?���Z��ۺ5���oxz�]
�Z��h��ݰ�y.-��[S�Qf�˄ ���m���&�w�����=�g'��::�1��}����j�/��#1|��z�+�4���������U�V�pbڐ�N��C C�P�N;�{H�ߝ$�Г��a:�_�\يC�e����#�A���E_��TF�m���&@�����FQ�<��2�ۓ�r7�� ���C�9+�`R��>C�$CWѡvny���9�
�\j�
�:�쵸�U��"���ȷ�^�J3�K*uK���"LE!�	��ʬ����ߧ�]B+v�V�R#�*�x8��J�UiP�7�7�S7-��Ւ�/��cے�����n���������|泮'@�j5�|P~^�B4��Rik���#�O����kc�>zJbc�	��ع���I��]��c=2��V���W�dS��,F�/�D�����r9�h���@�h����M� �p5�kt�S�0d�C���Q�~;P��d��Zᩳ�e��V�5L�y-�j����|�I|��/+}�3�V�A��"���>�|���P�[�����N�[Y�;�'��ª�m�n���'�dU���n�CѯM������~�D,�<�����H㛱(�ͦ	M�,9��b����	;���}@�>���Pk�>�=��xv=�p�7J'�����m{R�����x/s�tŴ����9|s�y�݅����x� |�vn�f��ȅ��}��R��ߤ˟z�X~�7���Fi��$�Q�Ή����ެ����\{���X�T%|�s�����:<i�E����=�*�b�]�Y%IsE)�F?��0�:Щ�jg�{�j� �g&^xU��>�]�u�edz6�~��e��W�����L�>l����'f1��S)^Ecf�87N�uj�m�Ǭ~�Ŷ3;��X��V*�4e�b�gDL`���\���-�1��}�骂UI=e�;�d�(�=>`�J�:��5K9�<����׵9R�y�5잀">��4׷�#�[zg����x4+"���W����;f�R����T�8wk����}��J��r�{��< {7�>�������xLऄEmZ�����X��l�ŎB���7a��?���ւ3ot���ql�f,�����7�ޖ\MQ�O2�f MPCa� v�d`}g$� /M�\�4�rAc1��S�����e4w�a1s�2RxÄq�5aB3x� �5��SZ��������:�,��-8����
~�,�����޸M+ӌ
7��?;�7��(U_�/ے�7��g�^�i�r���%SNB�>�;��S�������������ѝo^$/�U[����i��W��q͉�� �$��'��F���U�ƣ�O�#��H�Aw� ���#i:�c�@��c'8�0S�@Z�d����Z쬗,�^�� �T�K���q5P��e��u�����r�)�~��|%@b}�ڇ,�j��4������|�5"���)Ӎ�c_��:�/5�VttxF�nQ����j��9r��Ifk��������e�[
S���j���6SԻŀķ�+�8H���
�ha�|x�ck�V�~���'�O�DV��x.b/ŏ�|��ߗ����Չ2��d�>vwL�p��2e�U������LP#:��)*9G���O������_��tAsR�S����!ۅs�|�[��aWBd���C'L�i�Dt��'M)Q7c������
ݩ���:�����7��AvE��ō��߿zu]D5����c8���w������=?�ņU�vƽ����G����~L`C#��ͤأ�$_��6�*�EIy` ��z�yc:X���;���li��0����=�rũ��U6�=�O#v��k+<8��y���Z���E�F9F�j>]���\<̊�s��cc ��٪�����W�*̠:�������Jr�vr���Qd��(��\���<������^�U�LSV�����^��X��%x6�ҧ��N����8g~���Y:T:�KF���)f��S ��Y�H�R�\�Mw���	&�e#��<�;� �|5��J*�{]�?Q��=Ô�5d��vLc��T���Z�ۇe�ދ��^�4nj���~������=���Ƈ�.V��Dt�`� 1NJ	�3�-�wxE�1o�}��0�q���[񥥤J����X������F,|���g:]I��~od�uB�a}����L=fuG� �<$��-�-�Q�&�1|QG����@J�^���݃�&Q��t�����b��� �\��8�6/�������V��3g��.�o�g>���/qס>|�&���������j6��}h��	��:&ks�U m���n~��(�n�y&M��l��Mcc0FUQ�0�ܥ��,��҈S�Z��p ���g٬w}wr��>Ol�&���D��#lq��nO>Ǉ�+��fiЕ�Ѯ�Ӏb^�.��N�ٌ�pz���{8���,tNtA��Hes�O���̆���".�f�my���Wтvn?��&�+�3�I���{M��Imb8,͕�q��Qyi!c{k!��0�����Cl,׾����� ��7��gz�*h��d��3�d �`
�V7����lE��:R'.�w����!/��H��-wl��G�VZW�S���eX��{vf(n�'e����M錴xӧ��k�3[b)Yʛ�¼��Nfr� �����+�q,T�%0���X.Xѯ<��bø����×�Y=!�%�nnMe:7aJBn7���	�E�G�k[AU���k�|�=��c��z<TQ77R�a�&���hAĻ��<Ž�6 ��*��-F0p�y��մp�7���I�B�����Pe���Y���0T��k�y����x��sT9�S���s�M��Z���RL�p��&9�{AI��MP?Wۜ?ߨX��؎�q�׌��kQ�J�߹e�'a����3��/�H�!-�i%fmB����*�ޚzY8A�l�w�ӕ�,�H+_��׌U���ڼ�Χ�3<tS��O��z^3��"�J^K�dt���걀��X�R?���}��
��m�ri}Q{sbᗮ:�����N%����d�]�!r�*i-l�+�.�>|W+k�|�w��l���y�ߙVF&���s��Y����>f�-2-��m���=.[N��4�=M��D�Ҡ���5�������=��?���&���Bu��z&���$���i�I���I2������>�|�(_5M��ç P�%���u�W��n�kSXi��BeZ�)��'F�3I�،N#�̠ǀ��$\~0���ss�g��n�u����^ P|�:[h��R(�3�S+������w��)�j=(�H�݃"�2ߎv!V3�W8+�d&�3�WۉEyOs)	�F8�VkU��nL�X12.�S���B'f�[;���u$bF��]	�X�Qӄ��9������6u�W��(�Ѓ��U�G�"v�����Ř$Y``		/o���p��-���w?��sk�W�aQ�,��#a玁�~>*�����M�uX#�~P+������I��N��$@.�_��=�їQ;��=V��k}�\/gG�Y"}"b�k���H�N�7��o��k���ؾ���Vi�����\��S��pS� U��B7f�}�R|%���|��Q�Ø�����(��xT_`9��T��:�n��u��k[�( �8����J'�u��#�� ЫgKg���jˊ�3��������@�F6u�>bP-E��������F���F^-�c5ϻ���/�6*jn��^�y^2�U�����LXH,��Re��#RWy��f��"���;�,�pKJ�W�GH�%!�u���P�Ny��!�Glq
��� <����@�J>�����+�3�HV����t��Fz"����{��4����?֖(�~2�JU����^�C�ՙ�w�,I�19��g��\��K��l�1�1�g
�,+��f,�O_���'��ԣ�|3u���ђF�1V���0�~�v��U���R�m푀9�ͮ�x��ƌ��4K������F�������Ҥ��/��Wҷ)I�G�XO�ޚ�]%���p����p�ȅެ���p�����.ů�	<yb�g�J�pր2A����A�uP�Q l�]{�8�A�Z�㸜yn�#��z���+��YtM"�[^*�������y�h�m,kc1.��Yh�� 7����y7�,,\\ؠ��NYz��mߟ;��0^i�3S����IwIQ;À����QD�3%Z��em�>'�$�"���;����H&/�j��Y!霩�[b��u��\z��ע��I�s��g,v�Z�u�Zi��B�b�:�RS��s��H�
p�F	���7��"�K��r6��~Cv:`�S�����tx�P���\��Wlm����w��舠v# �ꑆ����c���'��"��R]�Տ�v���I����b��[&i��	��q;��o�45t?ܫ�V�,��*�N�c�p�$�n�.��Han�x=
]�9�����Y�
�<I2�����@/g~�%�&�HWh�X�>{�����"&2bSгm4�G�>���h�v}��,�}��u�iH�n�w&����j�L�1=UyS��P��h����E��o�|f�F+}��Q3N�6�#���gwRsE^��~K���{"�<�Q�Ɵ(#���$)�����/o)������_�i�[��z3�6	<�H>y�mu�{��T���8sc�M-R:��@�������0�OɼOm��ᢽI���~��6׿e����_}$�M�B�Q���ĕ�.���w�{�fQ����?G���{diNT����8[�@��WU�҇�G�/�4�	���뾠S��X��#u��L�b�*Iz��l���M�J@�|;���îIA�6l?|?`tL��v+�7�k��y�]o�
ׯ�q��Zh_�Si����#'�e������ϻ��W'�� LTq¶��ͅ��Z�T��9�W���z��{#i�q�r�>��O�/���D�z�T�G=oI��p�K�m�'f�9څx�[u�ݾ@1JxRg$C��V~��>�~�U�3:v������h&� �!�ݝ	=<�^�l�R��`��앳V+�9�W��ಸZ�K��p�/-l��F�<����p�W�P����m���t<���1�k��&$Fq,�	d?9���t;**�xz�B�-�پ�h��"65�oސG�T���+�����R�~��с���ٽ�:���Y��\�N�^�߉�"d����KT⸫T�⫌l���_UI3�}-*s��::�7�W���(�A��9�(�;�Y�0�	����1;\s�q�����E��j�����5�g��)]�]�^�|��ҋ���|�z�R�Q�D��$�%�`h��cԜ��'�=, �J};���:دv�1iP�g"ԯQ��Z�����P��c�
�ά.�d�4���o�h`�ZSrӓ��_�����׸L,�D)P�"t��͸���>	zJ�f6 �~�������laXv�l�x��,.M�I�s�u�M��7MU��#���9�-���^w��HE�H���ҁ I%�ʖQ&���ğI�6.��cŎ����=�R��<��4����[�rQ��|-�AN�H?���z�Cئ�!+\��o��@r���L���h���Vb�O`3]���)��"��~L�����T��U�����+���J�h�Z
���^��.�$�@w�'i�ȵ!]��c��v�M�a�3�-�3E��{X�ni�˯๩����'����5�F2v��L��֜���O���ݏ�e�PS/ЩU��\gc17z��̐5�e�����q��m�B{����U}� =C����RH�{�����%r{�t��� 0b۩���B���Q��$,����[��Є9�yhS�#{�D^�>��M��<�o=����}��n�4g�V�Qh�9��~�k��;�z�.y�p��h�%nKŊ��Ew_W�x\�X�[ɂ��o��m�v���̞CE��$9����=�BR'|�M�R���)PEH�Gy�a�Ґ�m�]�;�p�$��q/��r��H��
�>=��G�i�&(M0 T��TvM��k�� ��t�5ktp�Lo�ŏ�fb����[=&��ya]��a
�I���v��V%�L���h��Y����^����f���'A;C�N�[����	@�k�n?Ζ{�܆l�(��nQq�Sj�6�+/P�$~l�K���	���>��v���C]_ ù��v�O[։��Q9���%
�{�3���C�o��j�������cW�7�z�} 9
�A��߀���qV����Ғr|s��rm)�-_D+��?���1i��y��t3��������{k5+�P��Bl��'���7��T�O�R�`;�q2�� >'�S�>����W�>�!n���{�s�ş�\ڹl"]`Q'�:��۷k6wW08im���q�z9h��Y���1�����I[c���ahV���4�ޥ��O6%�kҚv�W1
"d�.J�Zq� �p[�h$Dׂ��j4�؞��s���ŤfdH�5t4Q�w/�(J>d=x�W�J��	x Ђ�5�Q��lYL���JϽ<�䵺�佝�6��-gAE��D��������N���u�o��2g�-�vȅJ]���M�O-�P6�q�9u�4�(
W1�D�;�����ߡ�� Z\��������r���q9�������[y�P��F��̯����t��#�ˀ�KF+��ѳ����O�ٱpM��dyiuT��{�����oN�^@
�0��;�7r!fs���B�GG,M��6Ɗ�YN}m[�.�W���jJY�1&�92aR�<�o5��0/r]�|9Ǒ�6c��ivFj�Tˢqʴ�F֏7�',	s�#�'ԍ�ź5��C�n0?��ӗ�썑y���c�"1�s�]�������/�� T���鰎7���FΥ�� ��ݠ���Jm�ҝIĦ~�e�<BO&E!,
^>ʅ)./�lEk�^;�d� ~�K����1h�l��g�"N�\�n�7b��c��z��sN�9�Gn�g
	iH����?�ʛC(&���Fa�����">����[k�;�4KŢn>�F��@5W6_���:�8��~�WR��I?n�1$1Td����5T�Z�]����`%��ㆥ�77���YzXr���Av���N��kU�?�������#�S��Q�^K\�ޡ�R��p�꒑���y���C78��m���kT�|3�tͯ����}��J�xy#}���h��%���~ܤ����yJA��F71��P,=�,��*����`�J����&#�jJ�q��}'zi�E�Am�۽�Ko�R��A���(���M�r�"d��� �UO%���m�+ݜ|�[B�u���v�uttW~���-�ᒨ[N��[����z��!Qv�0��}� �}};�Fn���KzAMXM�RHܭ�y��ͭG=���5���U>�+u�x<���K����y�����'�@���!>�$3+�h������h6��텠�jߥ�� �K�̃�%���:�xA-��\C���9�dD	�s�z{nb���?����*��oz�V:���ҙKGR�S���{�P��U��$����Y�f����"�Ӻ���s�A�����:�Hb�3��C��d�I���߉�}kb �(���H��*��  }�˥��ǻ�H����G��<(,�M��_�^��6}����y�pԁ��aT��C���O���{�J��V��_s8Fj�z�z��~�;�r�5�V.$m���5�~?ns|��\*d5OG4v��M��5�%�@t_��1�C)�k.P�x��!�K�Mމw���R�4ص(8��XC�=�D�y̹D�S*��[M��^� �*.Ś�)�ƿ1��W��gZ�}E!�&y���J�R�Q��C}O�ʉ��H�M|�<�����O`n�]~/�h�b&o+�oP� �����e&Pϝ� �j�c@YK��=$�)��k��c*��(H�,��W��k��{\�T_���һp��"�U|{�y����X�t,Q���5��G�84�)�8�:�tp-�����-�z� 7ڀ�oڈլ�/�I��9�(]�Jן'?���D�Ʀ�rr��*��2 b1���D'�0z��Bn��X�4��LY+zY�����M��{���
�λ�a}G���/�?����%�}}�s�;�)��W���qf�6�vɀ/=����'���\Ĩ=�Κ>8��UV�N�zŁ!�[���}8��F-�XeL�Xz��P��V�ܥ�FS���i���v��B��O�a[TB1Fz���y/q�+��wp���p�U&�ED!t����B��1��Խ��n՘ȣ�f�����F�,]��v��&�<_WvKه��G����n�y�/�r쓵x
0�3u������*��b??c\B�i�e9�SI"��ryV*�����Vz]ͽ1gŊ{p��Q����]i3:-�ms��9����sl�#dSLK�m��9�w�6�.T_��!؆qs�5���{^��f9�s���v�_l��}%��lA?��<����f�5e��C�p�����o�D������7�L��/X��+���t4�Z�����:�٪�����]������]��bLq������^}����P��xBCoD�⿊�QLk�+l�V��~�����3t h���-L��̡8�0޶�R�qn^�$ES�Y�ղʯ@�r������O�z�N�ӃQ�N������N�EAC�8������&圹���m=�@���ߨ��z���ẏ�_s|a���Ф���å�!�3�֋��x�v��f�^RP���;�K�j��LI�B����6�Q2��O7�����&�T͇�$�c��Q:��z0~b��Exc�,�z�����׏�w趻'�3fR%*�-]��3��Y.�d	���_�2�'��ꮩ��1{�[���1*x�'<'Q8d�@+�wt@/�����y���J�^��Q���>��Q�w��9y� �q�k]*�Nۊ�L�]Wer5<�ɦ�n4G��r4Q��_��+*4%�[�h�*���<|�KX�{u��a����|��]M\���u���[��/�\�L+������6TVsF�;PV#��ׇq+�Og�*F����h�d*Һd�¢�O��y[w!�%�Ƅ��"����r�d��K�?�R/�|��?�x��*\�q���:I��/x m��^Ypg�91:Xy�.x|P!3<|}���7�&�	!<�!��ퟻ��{��
/�T�H���}&�[����4�&���*p� l�s����$��ݛ���^d���`�Ŋ�,�Q&�@b�y���Wt�+����H�����E���iF�k��qL)/���;3׈�HC����-�� �
�~:�U0��7r�����&�O�H�ug�9L�>�j:Q��S0��o��Ve@���W:YQ:���(�xG��s5E�?�N�O���/�k�y���B��������5��s�t����^�S�N=�z>��!5��nf�2om�T�_l��g�ƃ�Lz�˷M0�NCI<-�L�T"\�r��K0Z��Kr��W�O��W�53*5#j���~E�@���-���lLHqv}\�U.	H��g�]&�U��M����A2�/5Z��NC���g�����08�����HB����rp@����
��W��3��U��++"����<e�*���9��˹EH���X���a��lӆdI� �V7FȞ�'����=�u�D����S[$�����f�>��	č�۝�}�9p�p�r��i��Gr{��Ա�'��s
��Xz^Ae����iEi�E���h��P}��/4�?��Ї�30Ҍ�m�ȴ[5�H��G������*��s	<����G^A�[b@Y�DY3Ҿ��}g�F_�N��Gy4fQ�^�І�W7��j?L�W��І�F~
:��(k>*W'��)�Q�Y��>���P��H� ��M����N乹4:#_�2�����8j/�͝u<:�n�`��Us'7C��7�@����ٹ�wOD�/�>W��k��"3=�mj� Z�!�N��NbA_�GM�Ћ-���1d����/����z����.�26�XԊ
���O�
]V������h%`T�2��?!$׵���<�z>��ˇy��m��X#@�y�O��A�Cu����R-Eiw���*`@3���L�\�w����n@��w��\Ԍ��/ԅ�,B�d��0�������>����0r3���%�˰�|�-x�6|Q�o�^��y �IgU��&7kS-i%Pï�[6q�l����xJ>t�R��+'��6��InV�������[�����|1��%.�M�޸(9s��%xs�V�GOrs Ւ5��`����*���e,��ra��jݣ�l���"\�0��c����{��=���Ķ�F��[�7,v�s���dk2�-��o.����yeۥ�bA�C��������^��Y�m���|2
:�=L�`uU�W��k.0��H�4���;��{` $=�M"�^��	?� ʕLڦHzE,��j��l�M�:��Zէf�:F�-'7�P�M��Ҵ�B4wNT|3 ���=A�M�S��N��"|Rv
�)�(y47���{d^@e(j��h�C���5������c2�%*���k�F9|�7�����e��_y%f���^�1a���b��ɽ[���nk�ϋy�&I����[��w�����.�Tpf�|���g�6�oٯf�K���(7�S�d��dX��g�{` ]��S��i����VfT[��&]��F�arS��R6!�����Sa�?Ǆ��G�"�֠�}'_��
�Ţ.�@�(̓��bW&Ԛ���}��1��x��N��ʉ�-1L�6?,�� 4�禠5\?��Xs<��^�E���w���=I��N��ۿvi�ߪ�q��6~��!@�f�l��-S���{���p����c-R7#����[����RE����{��mu��ݝ{Ҝ��-
�җz:��ͥg^.��w[LǱ��g/�r�0G_���{�Z�#���v?��@�=G�y!ɔ���7�r�ӿ2&=�_��x�W�.��iS.��<�C�6az���� 7��A��\���љW+��`�Pk����Ӭ1���������#=�v�.�J��:H=�ʎ�n��>�K�5dvyڰ�;�ZjG}�b�~�������Bm���>uB��$�� ��YՌ\��R�5�S��=�A�	�jT������q����e�̨_}j���oWƚ���Δ94�\�:�1ΤUY(4S������2��s2VRa#��~UD����4`3Ռ�/�E���\٩gt��c!�///���V��G1��V�?1V�hɁ�f�5��F����Ƀ���� �I������:��X�zb�"�]��?U<�=�Xb��t�<`��Ll�� =����wF�[G?��L�Z���$Qы�-�ע:��`�قd�g9,<%?��O�*��B��Z�6�/iXH�W?���Y�X}�Ғ�C�<-���}�X y������촩oj�5���ݕ~��-�9Q�6ݐ]�8��;���/LH@4t��-�3��U?PK����f�Qpt^@�8�@���������<���/�T!��zN�"9���𨚧]��F��  �N�P����0���Vڌ��\�A�y��)��r���$� 7�iD��/��)�m��������i?.��>�k�/w�\�Q۰م���{�\y(������ƒ�S�b�qǮ�z[_VI�dDO�cL�<�d`^S��g�}	o%ƕ�����(]�]n�ڈ
J��r�7�h�T���U(_v�=I�|��r�Ċ�f_�E�j�B���Q��x�},���X�A����褝�]�*)=����%z��mwp2�|<��a~ǩ�=��&U��z���i�����@R�>alϞX���$�!h�\��:�6w ��!�lC����r�5�۸�Qt�P��¯�#%7�g�]�0�q���[#��RI�' �,�����b>k��	�YO��z\ ��AxO��D%T�J�޹(����Q�c����{��ާ��L�G�YQ�>�;�f-�9 �A���/qZ9]X��*�����64�f���up�0!��7��m�\�\|s|~�9/ϼ��.��u:B�,f��K����	y�Ʉ�ƶ��_���Y~C�Mk������LLW'3�y3N�H�����t~;���-։q=��Y9��r��ß�%9F�x�ziI���m�I�J�/�Z�eň����.�vl���l�S�#����K�4 ��V�fD=" ��Y�s�m��o�.���lQ�kh�h[�������[XHH67��.�����MY�Nmo���b7�k��d*��B9�/�e�Z�� -�I�6�~�F�@���*���<�����U{m�묑����p=��
�y� 9ͥk���e)>�����XHB4ύ���c9��Q\.m=���y�[�?������-��6l������c�=�+��ߜ0q�
�~�1����i�9���BQ쩲=\��JRZ����9W���#��8S�@Bop�F���wb�Ͻ �߆�|Cf�d��ͨ����?�p$�ĶPEE��~G�F�$�vą	����tB*C�h�c-�����9ޱIf,	��9Mŝ�9�M�@�`�c7�yy��D˛�� a@���~�*à���F��~�S�6�Y��*�c�Re$l�l�����Zc�ېq|ռг������J���k�h���չ�n��z�0��(����Ot����,+9?��L�J>��"�?E�l��[$_��$���o��}-��j����I�?�3~�;�X'ᦼ)D��R|���J1��6Z1���-��c��p��Wt����g/�Nܿ�s�fA�ymn������������Ya��Y�n.(�{�Q�cI��}^���)�C�Ϗ���}( �\�6��A���� ���Y�zն ^Wk��ޭ�m�rU�n�E���P�>l��RO%6�m�"mjAJ��|�W]V��	��K��%9iO�Ji%���6z�J�X#�>-��<TK��Ph+���T`*�Jn�>!@==2�f��O���25��}+�<�����*#�&��I3�ܶ��5�D72.+ը�}�@ң�G ��W1�;� �[3���,	�t?�f���#��H
T��ꢞ����a`b�rsL0�����/ƌM���+���Z����÷�N��$@2Y�����@�$r���ά@�_�pm/�?ua��b)�����\Վ�0�Ko� ^�0}�����ߞV�0�����L��Jl3{�q08o�T��@WY:���ώ,�P�Z�S����P4Iط�D�y@;�V�0s��W�� LZ۟��Ě��t��'��i }˧Q���� �s���/+if�����S-h�ل�
�l��~N��Z\ʮ���>>�N���~��յ"'�éscE�l�q?�!�g)
d�0�v�\u�*��=%G��
�*�����a�]⩟i�Aϗ��	�{�&����_��?m��,�WS�D�z�A��}j9�P����˨,P< M��� �����z+�����6vG��X����[B�e���׈�9԰��2tT�X����.��uo1b�Y�j����|@�i¯��)��?�A�s'��6*W�0�&e�Y��n��� ݽ����C�[�+�8jƞ�����<W�[����S���� F�O���#��Qǣ�����&�%N�K�jv=��B�%�9y��-O���_����:�4��{�xn�E�%���X�m���G�x���z��r���W��xE/\1��+���/Q�C�w�{q�
;�����&���+���S[<�Oao��Rc:�T���;6Yb��"Ȓ)M�#w������W�5Ӥc�2���a�Ú���aQ�*�H�%D�"
҅H�ޤJ���H�w����;��E � ɷ��s���s���a0Yٳך5��;�f?������ I,� ���������w�~oT����(��,B�7 
<<��7�}AHaWX��!��~��P܇�b]4�U��~F�����%|P�<�r0yg\�@���g��z���Ϋd��B���	���[Dw(aG��k� ;�[�� ;����;f9��"줅�E��q_Sv��t�J]d<� �c�v��ee�at�/��:К�V��Әi)�Gsr�"��E�K���ne���X���5�}��o�H����v�zŏ���>SL�JY�O�˿� gF���+����쁁��A׉�^�8%���\`����?��X�^汫mG�9��	{oN
��W�N��u��)�0��@�������+{b*1caX��m+�_�qem_�����G��T᧾"�.ȧL�rX8�T�;�hD1�ظE�;�s�К��Q������Q��v�����[��h=�)�w�kn�H���'z�F���k�� ;�<�����S�C$��z�w���('7IU����lk�����V)`"���]"�7V���>�pV�<��J��4��+~���i�L�,�%�S���}{˦�wEZf��ψウ�� �x��$��V]��VrĖƒ�G�a�@����N����������o�KM���c$�ޯ.X"WE��p5���e3ܝ~!|NH��=T:�3�`%���G���0�H�>�_���Uƙ�0�R��3?:U	3H���̪�a\�� �eJ���p�h<���	/�B������ĵ$^�>h\"����1Q	,���Ą���pۀ�.��4���?g����r��5�Z̷�u�><����y�|���
0��td����;��������B��c���'��qT��M������xΖ���uC�h�|����=th�@��f3�ڞￅ�k�՜y����ܭa���%0��� y�(Q�'���p��	e�Uq�0;T�yٟ>U��ڡ�;tk�W�3V2Ҩ4�OKkz�j���}��ҧ/�������O(wK�I��:^x��)W����RlCV��f-����m��/��@|��YYp��|H<!T*��4� ��G0��0듰?�E��W^~�I*��P�G,A���h�W��̘�7������ݲ�`�1h�'�?ӫ �3������Aћ`B�Q���̌����$�&��N��+1�����y�U9,"JC8�nZ������3]I��2��Gy�}'�P*>��.&���At;�K7�C�7�/�-=m/?��џ��U*LPCD�3?/Y�9���2�˰�PI�{{����~Ӡ&��OK�.�����b�D[�a_�vV
���@
����PN+�� hV�ڬ3�e`��0��:�
�x� U��$l���3l�$�D��<cr6�G<�X	?�nZm����-/@De5�����Hթ��� �R�d�U�*gr�Ȁ����Uc���W�J�7�A<��l����I�TW:HF��m*h!��V�cK[l��2yf�j�S09z �n)�)q�2E%V��M���gO�~��$5�:��
��$@�vV�򃗫�;o,���&w�_�
�p[�6<��m�Þ���;�Z[�B
9�aR���޾A��)�KY�������I3Zp,�K.VWP�j�*�$_̥{=�F��	�V����h�:azɒڒ7\In���az�rj��1�����~�ȇ���,b�:��y���������oi��u��t�^k���������U^��S�~y�D)�`��Ȯ�]��&r�z�' �=�'L΢gC�b�����ϡ
pB2v��x��NQ���)�DJd%U��\�~�%�5��t�t��L�+t7�$�^C�ss�[�`�L-���f$�DB6�����/Shu�? �Ge�T
�V&-�> y7f��Ġ/��j�N�h.�WZ��� ��/�B��F'����뎊�Tuuz��N֌,u�Ŏj~al����VQ�G�[�,�(%��'��\����niQ(��L�`C7폾�d{-LA��CS��[\q�B��i(�bq�!�g1l$�F1� ?ԽA�y�hK��E�Xf�y�y��&&Ks:��Z�>�  � ����=�$�b%ݾ�@�]�8� Zd//l����i���A��FV�^�����8��4�2��Ɔ��0,��f�-h'G��A8/����"���	&d��"4����E[@t1�U�a�������!� ����;��_fn�rNy+i����DF��/����:�ʿof��,&Z��i�J��R�ߡ��|��y�_����=��F;*��$͡��ӃҝHF��B<�l��}7ל�\Z�V?����l~r�V�Ň�]�t�U{˅�<��M.��[�,XgO����JR�˄�w�;rMx-y�&��y��R+�\j��D�f�.��nvH^mR�������b洕&����r��ѭ�RV��U�[�'@��w�� D�xWT҉��R�ԡ��/VS	U�p�P8���ӧ����z�z�0
��P*W�l@��v��_+5�3ƭ�w�z�mNz[4��t��ݩ1o8�ͷ���'.�.���@ٺZ�n I��wS���t��Jb�.�.�J��05�u*��O؀}���� �
��f�]�.�ܵB�錥bÙ�=u��L��OA�����Ќ]Ӑ�Լ��vw�ju�D��ǈ�Q�gS�\�?R �Ly'
����K�e�o����n��w�[n05�P&l4�P��{��<@�י9�UïJ���x8����"���G��|H�r���~٢�,��Zc��z�����oer\��6�5�m�]y���ɛ�ia�D1'3'�%\�%�DI`(9�I_ɡ��| �P�8���B�;d�jM���W,m�_ �$�8��ϸ�l<�UH����W�{�K�qx�wL���j��s��
G��K��؎�>P�s ��+ ]�T��fǐ.�`��2���
�"�.B� �����0��Ŋ}���o|�L��OB��&U�1�66�t���1�pkA��f(��<����ƶٻה�Q�ܛ �l U��B�ӷ0���N3"ҥ?J�)W���C�ݰ̓����8a"�Wz�	V��$l�S. ӧ���lJ�NwRB��:�������r�e����n�GDֿ���O3HY��<	M�6q� ݳ�`��D�◆*�ZH��"󽪔����n��vZvǵ�!�h�b��"Q	�~���m)W~��B���,~En�%��{x�,S�>bv�E0��kn'u�ڐ�"���Ц��u~�V�>;|�:�I�R�a|����a��$Za�Ohe�ŔK��,�i��;yp�z
�\ϓ^�gL�[Kw��m\�k�}�f<(�����z�-q�j��KL.7N\���1���Mg,�J:�#�}���^��:o�u���Y#��3G��;���W}'ޅk٩l�#G�aLo_K_�G�,�"L�ɲۓa�yuZ��#b�L�hMu���15l��N-�� o �%�+n��'�#�V��5����:)���ʿg�-�S�u���\[��o*6�k�"v��3��n�7?S:�'�JK�y��mp��5��h�������)���C�(�~Ť��u��=(7���g��T���͘�5�7�H�CA��0��>q��oT�Hr:���o��d��ؽտM�$����a�1"[���V׃�� }�?��PVvr�F���c�D���Գ�4;L@��A�EP��#�_�'Fu9�]�K�����w�(1%u�<��ٚ� Y�԰;-Ab/8w��
8�2(6}�tq�k�?�u���a��b�E-�x-�E���ӯvP�We������j6C8�g<��;ƅBM��-����x���ϭ~���������4r`.f?KN!{���`�� ���.��XFe�w�|v-���l�ϣ��� �c��פ~��-C^uC����q����L�S� ��7�s�B����*H�O�z�����nPg#������"����l8c��u�LW�L�����ܻ9�԰�԰Ϳ�G�K�R�M�����Ņ��q��$D�%�O�\�D��� %i�d4oJ��|��rL�@����o��k%�L� R ��I�@$�����`n�e�klg'�$2�X��Vcj��3D	y�,cO=s����HXyAQ3���.�*���v������7��RL������ב�+9��Y��D�U%����Dk�3��h���D���-�Ki�mm^��O��w���eΥG�	
<k:����Oa�L$olia�x[!Ò%��X���vq��Ԝ�[�h ��[�̟���c�Ŋ[�
�M�)a{��@�d`L(5�G�*0�g׺����>��j���� �?�z.'��%o�V�9������6Ȗ���W�t��8L�K;���Y��*��>(���d�j�d|P����s�O�t�0����8ӫ��	�d���{�o�K���O��X��r6O|��l����m]2�2m���ǿG�������S�^̣pK�#P�E5���wX�>��m��R(�������ݚ:�>Q{l�or�O��Z�14&AlW�Om.�=rB6��ye��_��?�޳�qrJ�?0�dR���F�=pK>��	Y��#u��D�ӘP,*�{��qV{'�+�0ɐ7N�t�F���)@.ݳB�c�9j�Z�]�fIqH����+b�o*�$���A�l�{��I%4�4�^�`����o�h���e�nq�(��$����IX�a"*;$���􏮸�1憺�ƶCdA��~׾�P�ك�o::��\��
o�ǜ�@��2L/��N<j૨�r��Zvr������;-򒅃���;����E�ëi!\�YrR�k,���0n�nl��5)n.@� տKsi�����J�7�o��\���tA�A ������T�	�PO·��{��/�$2�W��=�GL�	4��c�L��xe����_��;,N�g�l�`�˄�{ ���;� �p��B�����; � ��S�	�:Pr�W������m�o'�3>�IF��`�u1~]5��X�s%�Y�k>���]хsN�gNωi��|�G ��ri���?Iy��0�� �E�v�X`ۺ�l1	��)�B�"D���HE���L��sR�KO@�pPbx�4@p�X���r6�as��f�05H3i�;�ˮ�?U�_��9�BICK�A 0B���������R���-ǵ��ص�u�d[wzK��!���seM��s�����M�����_Q��|=�O�2��{J�}��:%�%ה����yS�B2�&�HdleO�	�f���!��>Ha�21@r+���{��]wq7RV���u��#�+V�p�n��;3�m_����o]w��L�1�sjgi���v���CG������0%��}kF��I�#ub��0�AgY��4����Cb��x+[Ϙ�P��Q�R��}&�@�rߗf���P�Dӆc�~�k�p���ov��Y��m�-X�>#&���F?#�Ӭ��ڤ�#�]�)�����TԔ���nwE\˟K��V���^4��|ګ'��ΐ��ځ�#�χ.&c����!�V�&�$�^��j&����֭���k��TNY�
���1�[o*�ɖ��{�3}������8/�����*�U�x?h��`G�hx��J��D�� �44������qe��b��>��`!�E!�3xr�4�m�J�ǟ��I�ɗ��k������fC`�~c�ͤ��l�d���}��w�&2"�_�8���C���XV��h@ؐ����.%c�zP��e�V�/���̮T��ч"�3�)8Z(U� @�O��5	 �c���$�o-��6��l����*�?�W4b�ʞi�))3>'4�t���gJk��?�i��j)�̗��{�$�Vk��C+ �w&���b����sMidƐS�q�r���z.wP7:��mpz��ǲ2��1 �J!q!
.�>'�`^���1I'��V�w8I憮�6�K�4��TH�r(-!��#�W���A,��d�~������`#���V���@ځ���`�T��i,�{ƳbG����J*+�J�����1
���\��P.\��#,�G�F��{E� ��9�4#Fc4E7�:� ����~'�a����פ�n�N�׈3bu߂�^�t�}�(1�O��Wj��k��O|���Wu��3
7����J�d����Q�0����/�m��Z�6�)���eh��W�_�;V��ë/�����A�E/���0kw���D�;$eȧ��\���L�ߡ/Uz�[��.Ҍ�yI�b��1[���u�MX�����)���Zf��R����gl������`�43��.w�n�?��}.�1�\%4:� k�S��Frv��[�}���]�����Ssm�q�����_�ڠ�)�jx��� � Nu���5�t]Yaͣ�s_P���أ$���OV���~��zߍ)OZ�&\<|���b� �q��qú蕋.TN3���:��'�9yB��_%�ri����!�U��	�͈G���Xe��Pzvq?�H̽��~c��Kſ�<O�����ܓ@⡲�t�p�H�
$p���h�zf:�1i�D�?�W���+�}IJg�X[6�]$�ro��_��#N��K��&�l�=w� Q�-�5���F��/gl��6�F�s��#$����Op���&Gd.
�{��������#޳�@f�����n�i�R$Ӑz�����4��#�1_4�6w�6����;6�9��S�Gm{��� e�5ӏ�Z��ޛoL�J�=��ه;ۣW?X��U����n�{���ǧ�>U�,�����K_��d����	�X5/�WI
.��kT�x��p��-7)�E���;��m�����7��D�μ�3��'2�ڄ�"w��{{����C#�K����y��#��E���IA}$R��G�Y��F�&L�c�n>�-;>>��0�=X+O���_�ߥ;F�S�*f�%;ߙj�2��CU�}�h��C������ۅllǙ�u�F6�<���:�hR[����氻��,'�Ӹ��'7!o'����VV�bb�HU�N��ҳ�b��B�������	�yC�rO��&�Y+'M�"�Z-1�H�Q���[�MO5�#���WqV�w+�U��Bߠ)7�R�W`��m
�j��m8=O��Rl͌��K�,����.���v�iyI%
]<U���H|�u��@��@�ԥ�сʴ��:v<Ak)i<���C'��/0�J肜qd�n6X�B'qC<r����U*v�N�ʡoWb3�C������acV7��~gy]�[D��O���&$�G�g���
@&w[���ҋ�Չ�o��O �'�����z��/�����OE����*�^:��)��P^�|��Wϝ³�*N��8�FO�X�48��k�������}��Ǡ���j��Vk@���U�x1�~ �w���rp���h�#��\�r���K��O���	fF6��" }4���[y����T���w��3��"n^��{v�$����㰑 �߷��9x���Z��ׄ9�26��yy��B���g�o��nq�K��{w<�ֹ�wMm�6�=�!|��ޘGܗ-��L���
f�c�US0�q[יJ�@�l9p�B��鼮+��ty��mtX��ˤ1q�c	�&�����n�ꁆ�j��B��ZULp���F�7��)��Ұ�,�{���
����Ņ�l�â�q��=�;EͧE��l<�f}a���%	��&����+��J(�̃��)���WCc������vֵ�4u��k@촖��íѱ�~��QY�j=�ZG�b�wWLM}�J�q��ڿ@E�x6P�j|�wP-����q��\�<�s��v�����g��O�L���r�����-�o8��,ͷB��&�DﻷhBF�I��N�4Զ.�V�rY�����;��cJtG��P�l����^�D�[�ѿ)�R4s;���e���O܍��T�q5����k�����|V��f�=�Gʻ9��F�G��ƌ�
�W���>.��Һ�5�H��H���cߠ`��gJ�wxɫ���8s����v�1�0��;4a�F{B������S.��e���Mﾐ�i�׭�� �E/�b]��f�C�/n��SK�@�;�l<�i5h��[�@T.�y	oІZ,�7=�8�'��tcB���q�u��8�o�NO�UcV棁H/m��w>����*����i������1᫹i��T5I%�:SF�P���� �6����1��������<�d2^phh�����t�a�������l���K�d5О��b�^��	�s::��z9��鄃-��<��~�׮��i��U��`��U���~rͭJ�ٽ#�Y!K���3һUIn2���g�wNl�K7�c~u�jí��K�X��N�Ӵ3U/����kp__����d��_�j��3nzm-����9f^uKO�@��f#'P���S�!]F]d3LZ��IQi� [)jSn�@��B����0o�\K�k�Ȫ魦Ja'Xݜ�h�8��%��8�XnE��n���Ă	{����S>]�;��ѐ���.G���	����6c��G;f���6��c{���/�����ӑ�z��h7e��϶{�[.�ӱ��2�tmf�'ӲT�yb�aN(��"���,��#z�nM�yTm���`��_ߕ���k&�{+�^ϵ݃�}�.sr��\�R�����-		Q������4�C/=�g�.Ř�H=۟?W{P�@u�lk������L�E�f���*���B��N^粺� ��n�,K�=**7.?�sw.�h�y�P<Gw��y�}�%��B=�g���
���2z��o<���`n롰W�@Ч#�-���o�3��<!jp.��U��c/�6E�9Ϝ�U3q�cݾO	����&�8��ړݝ�㆖��� ��r.���6\o�Z�k�X1*GV�Pi�4��p䧓2��a��TK�~�b��@�苐Ǔ����\��٣�A6�7�]�$׷���+:Ӂ���ת�O���N�݆�4&����<�<���o�rv/Gɮ%��������aE��b�p}eO-�H�1�s�~���0&��J�۸R,�6���í��6�jUNj��ݛ��ձ�gJ���V,�	<��ɫc���^�UX�C|�>~��W9}R��9ioy�>�k�%��?l�;��p:���
5�`,�#S
��8d` Z44Y�1�F���lwnm��O#bO~F"���j~�M�ob
[j럲��_�4"g �H�����Q�@�h{@��I�!đS�S4�gᾼ�(p�l9p�H�e؛\:���rS�r=�z�����[�[w�ԣ���B�7��=Vtf�g�t��L�-�O{u*r�� �nC8�n�b��҂yY��LCpy 2?bp�ݳ0��L��f{�LyޘR'�>�Yⴕ�������f/���p�|���[�Ê�Ƨ�A{{�;m��&��= b��vkN^�F�~DDC�g"�B����!	��n���.3K=����
X�8RX��˒[�VsI��P��Ja������j׷]��Y8�+��)r zΩ~ݧW�Y���>�Ҫev�ݔ�6���D7�ѻL������ޫ�����r�BD�49����UR�d�r�ᖊt�7�9 ��5�Nʩo46"R��ؔ�����+I�Q�UI#��FS�$k�.B���=����]��Ff�MY��h_�߄q=o�F�N'�5�I�Rxr�H1;���B?���J�y֧�Wi��<a|��v���0�0���i�Ӗ�un�5v��ih��	|��!0�6������ꪷ�)2�?��͒X���ƨ�Q$���ҧHI����O��Q�d4r��Ӗ�hhu�U�3,��O���8{u����FbI:�k�/��o�R�V"���s��)�?p/ě|Q jR4���ǰ�/=�2�aO�60G�?�8���"%f�]�v5pR� 3���N�'�k��foe2�L 1T��klc ���"��`Nj����HP �:��_�˱Mx�5/5��t��nm��R9��>~�"�q�f
>	�#C���T=��1hU�}�?]�;j��~�pr(k�2'a��D��k�[�iE�����wV�	�i�3���xZ����~2�`*ɮc܆>\\��F �HdC�f:�͎eU����}���v�I/3� �'����El�{�"����1�D���A��A�1���{�,C��
xܓ��9����	����nvku�lBQ�5Ck����a�[�t�]�G����6��n����p�qco���6lhK�;CM	�|��Ma�z�S[��<�3v��a�<�D�[���3:�c��x5Te���I�d0�*E�u���LyJ���S)�N!9�z~$�
s0թ�H�����-"P9ݯ�1]��s�`�p��7�z��IN�x�͌?q'
<E&�p.������_i،/���9 4	�<A`i�PE��k Kp�����n��Q0�,6����� b�b���"6!Ѡ^á���=��*���ٽ�<����1�\
QR��I�/���3�Y���ͫp�!i���'���߄�~:=�����}��40��E��T���\A�_�h����P��ᐉg�03���0�C�>��nU��8n��#D�����>R6X�uXcb��l�v����sD+g���9�;n�.�OI�q8�i-#i�Ļ7����kэ��7SPz@����̀���A08���2�JX#l9�
��d���%��v��nJ��UL���Rg=���|�m�����5�*ɕ�nQ�LY�D�F�d���-�p��C<��n��7�ɯ�iu%�<��K%�O��]j�ځ���`wu&g<������I�_#��Ӷ��L��TvE����˝b��?��u�����?�%�y40��k�R#�9�g��oV��@7�l9$#� ~���䯄�4����΅��8��#\��
�Q��S+�up�'!�o/܁�s'c�A+�Y��~��ۻ���'.�H�R=��������c?j�Ieq]JZi�t��S����n!��ES�l�2]���'��^0�Ԩ����PI��7�_�g����'�[�9b��f��|�b�z��ҡ��b{Ep��V������!�O�?�'�7V��������s�����?�*�,�ĳ1�!K���+���><��|o�'Τ���۳�}<�0"V�s���\�i����{$��a�}壘GO*k��f%/���8�iE^!�^�gYw�eU��I=��Z���������D��oߔ/�Ö�p�������1T#��FRLOeY��T��Q���o�ʱ���Bz�I+����~�E@��������dWŎ�B�5�i։."ą�����TB#�#�Ae��l���7Fx�5���Cצ�U!b6v�[�H'L��*SDr�� �����1�v��7Q>j7S��6���^��F>2%:�b�к�Z�×n�O�\�(8Q/�b��ψj��T
���n�}��X
������D���[j��)�6���h����J�_��WC���Tkm<��S*������%ht5{a�4������%������M6%e�!:�j��ӆy�>�ր2����/<r&'���'��>]��PZs�U}v���OQ�[���h�1�֢���[��_�
g���1��!��N����:��v�:�p����̌[�hgϪd��C��+�g����0���X�x/���wq{[�Z�و�n�\�9Ɉn��5���mu����+4�Ҩ��;]yJ�EA~�2�p�se�:7%�g�����{Pͬ���!���H4��Ր yY�'-D{h>����r��H��-֑i��Li_�Y۱��G�wz��T��nR��h+Y8ǷΞ�M���9x%��e�cy��Q�!�!���j���1�{�o.d̦��eF+XKힶ0�Q��_��5L��g]mMȅ5���,��`��հ��]�ggZNf���UE�jky{����7������b�V��}"�K��қL��AE��_��&����2�{�
�~�i���g�%�uk�r8t���[��/�ȫ���i�������`�O���U��22�����%-j�871>Dp_�E1�vܩ���[��-?�Sxn4�&h��<x��q���De�����
�&ϥch���yjߞN���s���~N�h��L�bw[�h�g�����kyc�e.UG���Y� p�c ����*:���Jz_�����nn��7��y��RW_�!ż�Ë�ղB��̚��^����o��|Q"q:���m�R� ��US�֞D�c.�٧yWK�9eB��V/]��$\�.�u�g���
�6�ȅ(�K�P��&��K8q��M�߳Z�ܞ��0h��2|=�!�L��%'��)��Y��_����4���?N�+��*�Z�N�0�h'�033;Q�\-%U��x���=鍅%�餱Yv:i\%��,:���#(Lƹ���rF����DI�;��4�!e�)��ې�`�0s ��=���+��gL��~�"�k.D"�����%z���#"d{��֯c�[ѯ-��yJ�p�Ӿ�^h2�ï#XzVtG�l5{����K���5ʚXKQ��H߼�ޑ&�����d�2c�7�!o�QNf�(x͙xFe���|��	ָ2�\��h5q�����[c���T�V�']o���Tߌ���_X�	��Yy3��SF[ǓǙ�%H8����Z�S�hJ���ЧK9����Jq>ݖ�X��{��;{�[�AZdX�2�и���V�h�KM![ϥ0R��*i),���N�y���_�NWV�Q���MȭBز��5D�5�2����G�ѐ�����n�ǝV�y���&�ޅ^<�����{c��n�ϋ�Q�T��]��^�36*$� �n�Z�VBR�uݓkw���q[����ve��������3]�NlC�>|����+y=W�*�Ɨ����ſ�#�y,3t�ñ3�[��.[.���h�$U8��ɲ�v�X)E���_7�N��r��}��8����Nv�K�6�� ���SQ������/Zͧ�s�ْ7�3⾞a~'w&+S�
��'�ȩ����s�fv��4-z�]yd�9*�X8h��Wݧ2΄pT��p��i�?r�D]W#� �{��8�af@<��W�p.(�j�-�i,��?����۹������''��2�� ��~��?9R���u���`�MF�R=��<u��@d�)tPL� p�Y�d�������W��$wV0}y��W ���$Qty�_����5�����&�+&㢚�t�A���A��^~��\t����v�%ǫ>%�v�軕�_/��8�i�~�IC /�Y\����ꏸ�xC�t���_AG���7h?�.|��X� �RX2��,1 `��k&k����q
�G�����pqC���x#�<}��s?Slz��ib�ɶ�����Q��Ƚ�3��\<R#�y�_vq�j�ֱb6*_�~JĐ�����,���s���x@��-�Y��X���&��oWv*��a����}��ࡗ��i�e�d��7Y��q���d���Q�<�o߼�o������F�r��^�n5�k!P��M6�sâ�w9�p/�Ӿ	3�ҧpm���4���^�&n{S�����[Q|ث� /����l@�L��u]Ux�hpu��Q��9��S)OD�ޡ��e�p^��`	���D�+M�"��Y��O$���� �ͺ�U�):q�-y�O��u����D��{�� ,?���$$T���Rp:qD���/C�@����|�����@��PӍ���G=*Z�oRt���eD���"����O7��YIF2��=�h�o^�#���\
=O��UGy�F��r�`$��c)).�k4L�N�jH	�:UQ�Z\��)tW�o{A�uu��z�0��b��=E[7>�,�(�<Sޝ�pI�J�u��{ޖ����v?/�L{��w��-����	������Nb���lhӴ�Y������D��Tf_>t���I=l�u5��J�r�%fl�½���T��ϯ
1t~_���B�k6'/���_��>��C�O>���|ض����oVu���aA��	}?�g�r�}d�qW!M]�|s��6�n�N[������@&� ��}���E���@�,�����~����--�'s]a���`�������(s�O���1qm�.n����z��0���!3�=���7��7#�9�T�|�;5���:THs����$�7��3}�u��D}��Jކd�lA�%3X*�ql�1�������3+�/5�+&8��N����d�,>a��':s���S��d�e�����z��C�:�:��`��\��(�s�
.��xE���#�����7̟\0d-�}�`YI����m���'�Γ�πfȨ��jK�^?[/Eu=���o��@�P��щ�C��(��d4>(8�����J,S慦�э5NP�|���0�c��w�-�h�E�����k�q\�I�$��h�>XL�๻P��b�0�E&��#����ڬ6dF)��8+܅�ڑ��T�3<�,�"ꗀ�~�D��Ч�<yt��E���_łk�_�Xq�M���sc�r��/U��ؖk��=��{t=U�fǃ�9��rj?�d联% ��Y0dg-r1'g	���������PH;RR���I�둯ё���"}���
�E�wf�� jo޹U�H�e�޾�|���qI��w�ɩ��M�>fLF�\M�}��/�}�A�-�V���g���C�Hd�i��T�k����|�}D�v�n�#k���Փ���}��I�ˌ��N.�����M��22°5 =�>����ٮ�Z�yH����kM�~��Ջa���A�;�0�n���騝�c�'�vи�dԟ�|$&��+���
��@��O�/艟��.��fi(E�s;į�`㟣f�X�C�.+CA�jC2_b
�tX��Ƿ΅Jf��a��SZ���b^���m?2X�ЏaZ�ǋ�2�05��M}A^�[*8���Z4Ƣ&z(m�Ir_豍�S���xkwW ��>J7,n0A�6�cK�BK���ƍix��!��s�ȣ()EC�Q��xR�眩�������b��F�������+�s�ˈQ5��l+T����1��~s"晕�22B��ͼWw(W�����[��A�nr+_"�r��ܠ�N,�''M%����U��#g�5���H+U|S��P������_âz�H��&tچg��ps4-u���.��L��S�����{�e�7tt�x�A���N����El�b�y��#~��Y�%ݘ��2����t��Z�ܕĜ��������}�~$�>�yZ��:g6��f@��g�\��S���9�8FȓR�_K��%u���8�H���6��}^�X�DR�}�>�?���6vS���U_�Z�D��5�7��&�b�?+������[�,�있PN���x�9&z�t����l(_B�2����J�ƢZ���_$RK��U0M��0;�н�,��_䙞���K�R�s^bM�M;v- qP��"/^A�En�U�y*���0��,cL�:����L|��<aZ���7���/����bQ��	�Pܳ���L�PՐyU��=���怯/���c�J�ɘ�w��r~X&DK�dHu��e����H!�����Aȏ�bE.du#�r���lۊ��Y�1�Ϸ;0����=�_R$�eu�5�ΰ��Ҡ2���x}�!�6�
��TqQ�+j����T\b#.�}�+���О��ϠCpt�!��e����M��S�ND~ί����:b�������햐���>��s�^,.�`�BtYFI���_~`ɯ��~����N"�m�̘(#��h/�~ka �������ؘ�^��_Rw�f��j=��%���L7�-T$�G7x�1ʞf�z��d���š�޳��O��J&�SO�]U�d�#O�I��d$�g�q⡍�{ ������U��DU�J 
j�XD��ZsI[�Jwފ�m����Z<�H���u��9�o{�Q�%N9[
� �<g�C2����~=�!C۷��rˋ�?v���~�;����䕀���ܞ��"�kd�����dQ����6 �d�ʏ������B����S���l���)Y�H�v�v��}wv6�j����ٖ�~<?�E�?�RF9s�k>'*�.<���圔���-�צt��[7��L����'�hY$H5���g��%��f_��gǥ�ₙhXפ�3)3�b�sVO���r�ޯ]؊�-��N���=56�L׭i!9s���PF���C�ќm�At���0�^2��ZO�El� ����`u�Eʌ��$/>[��M_Ա���yR�g y�������(��~-;��n�&z^ҁ�l��h-Z�R�r)��y.��0�b<ٴ�V��Y����V�w�dGVR�w�V�������Or�Z��B�9;��cڱm���D`��F'Saj��w�=f���6%�x�]�Z&���*�OD_��[o�/Ԧ���i����X�	����۴P�!u��+y�b�u<�/V�KތP��]�u��Q�����JL{lZ5�}ġ<�;)oi���J�b&��G��ŸVO��	͖���g�sAk��#�l ��1��k���TsN��=KY?*��c��
I�E)�p���x<����6��3��X�d�1����&�h��:�\,��Ge����))CE/j�󴋫Z�#����@�$|�͌�)����Y9NF�]A)l���ϳ�j%j��\�⾂t3,�_�V����7	iFH�F�ETd�����F�"�K�q�� !!%�hIa�� 
��@:r�F����ŏ���9�s�;�u�R>�Ub�f��ê����'��gJ�u�C�8	Zl�Z�m�iѝ:+��h�
o!�a.����k`!,�+?lGr�F�Zm��֝D��	�ǁy�T��S`����x��X�Qgm���/��V|��݉N�5�d�
=��Td�㞫RWx�[��F��6x�YS���?x�d�ި�wc�Me�+R��ՄO�Jhb�8Ốt�0��W�E��,$�퐧/�^p���|��sP)�sRcx^�`f���g�tFU�e/���q_���$�_���<	��Ậ�_�ڈz]�A؛&�Q���^7�1R�T�8Q����3�Z���ס�N謌.�׍���]~؂<S���0�@N�Yi�i�-9��H3}��%?W0q�s�(�T����`�z,r0����߾���K��������[��?��Q��q�QA�0$ړl�*˷R��)����%c�ћ������҃�Ӧ���u4��}u�Q�V�ٷ�L�ցaۻ�ap',7m���i��1g~�����L䭏�2E�Em�#��	�ʅ�ƫ�Í^T�蟝Ⱦ'��u/��u�N����Uf�����N '�O��S�:��X��/#6�A
��rd�d6`>Ȟ�����	��K}������g�E)!<U�\�M��;���;�x�]�+	��P�o�Id��ע����r�����.��d�}=���^?��� X�7���!�b��u13�HV��_tGIi����L,�uؽi��)6߸ݾ+�ݽ��xfq>��޹�rDN�d~u�N%�nY[�O��>�O��j[�H�85Bn��j�	��쫟k��{4[yѼ-��u=��{oz�R�iO'��Ǚ��\�������g����m�{���H�|�բ�\�v=1��-F�.)��Og�J�~����y&�nq����َ���������]���]��ot]��\z`�	�"�Țϙ�_���!�j���}1J�r�������פ��]���2�;Ft.�@�����Ö��$�Ѯ�r3���.=�a`�vH\�o�!p�-Ȏ|�;�3���2w��h����İ�����V��X������l������[��3����#̆��WӞ��R�$~b��q�Jre<E_��]-�Y�h�RN1]R��K$&�L�C��|�ޔ�s9��$EVL3`5���H=nQ⠱�ˈ��t(�t8�VX#��J4�Ķ��>5��~(�,Q~&��s��Z��&�8]�����L�kRom�)���e���O�TQl&������c�]���)f2��C�Xn����Jw��HC�V.�ҟ�����C��(2oTd!ٌ2ee�Ƚ �r1�U�Z��t���~��5?��U{��#eU�Tg��l� �TEe/(bv��~�g~����N)p�LO�,�Μ�e�L2�l���=����\ �$�w�������m���%-�=��,��L����0/�S%�� e��*�G�q8_f^��ǅ.�d���X� %�a�K�1[y�+;3_��a/�%ݼ[�5;����*7`vzZЦ�� @���+��+=o�.3~!�Ժ�� �G���[��� �=^����y~T�(`y,�=d�`E��1�-��-07[�^d R斫�;͐�.��.� -hU�������1��`jcnºe��r<�����nD$@�{�\�]�S��S��;o�ٟV��1"��L�;r��)�������u�c3�d�r�{�$�������TV���C	���n�����^�+�)w:�#ms��kz�;�2����4t����$�iS�5��R�g̓{��(�@����pF:�+4]2Ւ�/]�2ԧ�!X��I��N��k~SpMO)���ɿQ�(���`����C��]�t���J�2��y��G֪.�$��{I�	j�v=�:�<^�E�e�6��V��`ɿ���6�_}��`�* K9��4�E�ֿ#~ :H����C�n4P�[�+Vr���~k/>��.�~�Ӥ�r����&6� ��x�����r��]ZT��� L3S��I�O�K�����*��3��2�J>�ʋq��Ǔ/�s��j� ��>�^++�~}�x�Å襥8P�n�-gg�ujר*W8��h$5%&b益�C#�Im�����ġ�;�Ş�
3�������<���}���;�	H��D{<7��>��R��x�k){��Xv��mn��J.Z������_���+��(�����#;H��ߞ��6P�	,�m���9}�����90�
���M�$&?1���I���M��K8"���#�W��v��S�>�3��w�����Yz��+W�n�#�Wz��4f�J,K�Դi2��@��t�����|�ј������Y�n��3��ݶsf,��X������e��i�Y����X��o3-Й��})�S�Uv�zɂ���&�>CϹ��!���v}���f�����(�=MQ��M�b�dPN����bw��*M;����՛� �數~�?�{���7�����$Bi1��Wn��#�ٖ5�z+S膑�c�9�	Us�p����_��������gD����1w��=�=������u�'[`�ŭ�'W��"��ԁ�#�ݗb�.�}�͊��f��z�\L��k-�^�$>��sL	�q���S�H~E)���<ch�H��]?L��j�v.$�����h�����`�����he�h�Kϗ�-�	�^���ݷR% Kd�):P|
/�z<�6�f\k��2W��i�	��/�W�J�?�f�7w=5��cu����iHv/c�.A���*�q�Mߠ���Qؼ������t�ۻ�LH<�W֌!���֍�ʠ��(�FE�����hC$�������>���uUs�?�>�j�Z���i�̄X^���NPch���a��b�IC�j����ĩ�~�n/���j]�(5hw�t�����?���Cf{�c��N@ĢN�v��:�Lt����?%�BU
�p/�T�D����� ~H���}x�0��zm���]��i�m��#W��� D:�H����/�"*jc�7�ŵͤ�Q�|��]�$%�n�H_��v����X��������������_�x��n�X��D+7܀δ,��*U���A}����GF�<bN�k/��ItB�7w���egy�@͐�v�����m+�+�M�\!g�3ɷzn㓘�+%�zt`����4B��J�t�j6�fҨ�o�J�`��l�R%$j�컄Lԍ1ل�X������fL��z�X���?����1�
��c�7E`;+�ѵ� ��V*��`��M�],��S�[����.١���y�R�v)h��0�l�L���-����O��׶�n&]�����E��,قύ�������%)�A�\�_x:�F̈́�"����+bz�G�G��X�U��'X�KP4]p�G��OЙ�_T �S��:��:�Bj��0�ةM�?!�u��iI��!Odc	L��*��l{���q�v	8ch�
��73�>�4�����1�}���v�G�HIp���90�E�m/=���"�I;/��&^}�����*7/�6��Ch#�U�Ca7��q�DC���©<���i�]�֜d���Om�]�W�뽂�� Q�i�YӔ���I�d�<~z���sћ�tu ����@��fJ��c�i�H>	����q'O��[ځ�#���s���)]	/F X�XE����Nw"��Sj�)�@��*<KC�M�id���TyY�����&͊8*�5�6���7!'e�	u?0��ZY�J<�[�zz�UHN�cA�W:rn��;3�~L
/���0yӨ|�r!�3��oѴ�h��C���K�@i`kV��Qa#C��<���DZ��QN��9�C�x,�����@j�]�dWO����
*R�#�5�l��;��?�5Rl/V���3(tt�DڹS*ѼU�+YQ�(�5,�~�ICr"T�^�����&�Osd���15��&	Ī$�1!QG��Q��i�?PK   9l�X�o��  �  /   images/54b474af-19f8-4da8-b85c-ecb600c58ca3.png�q�PNG

   IHDR   c   Z   �N��   gAMA  ���a   	pHYs  �  ��o�d  0IDATx��i��ՙ�Ͻ}{�ٷ�,��Jܐ��ca��LUj���T��������2���ofR&�)��K�d�(����&(�"�
Mӷ�.=�������+Ц���C]��=�y�y��l�t�]����"�+ĸ��[b�رc�;��wG���fseee�T*���e����D�>����e|N�緄�^x���kY��������3����Mee���s���W���&��|Y��B��/��������y�9Ϙ����k��w�.��N�<ޓɤ�����R������"��g��s:�u^����l[[[����?>k֬�-Ztȷ����x����}������o��:�������ǜ����C�����\��|n���߹��'N��>�s�<�O��滟�knn��)~q?��L=��sM�3�w3��]8~];y�d|��/���?���<��c��^��_���׈�`���ټy�}~��A
�ooo�'�)��^&!��]8��}Ў��t:m�۷�}�O����b�A�C>w�$��^<�K�����|�D��}3o����UW��X}�*������~x�<p�y�q����_��׿���ы�u�@���W]]�]g0B�O�:e������I�1`���.�@t�O;�d����%��^1M�����Bs��%-����=�KR�;�0�3g��sໟ��z���.]z��y�>;+1�4���x��� �*��L�k|� �"i�w�+�=ЇT�T ���LĹ��g����_�~q�R��ڊ!�Kҭ1�0B��:T��<0��H:���cm ���h�-[��_��k�ظq�^x��z�ä
N�>m�d�ٳ��ڵ�B;:Y�����k�u#G�45�����ę�_�i�&���wA(��R�M�殿�z7h� #Vw�`\ ���O�_��o�Ý�Qc=z�!��٤���㣏>r�w�vG�1��xŔ~�vÆ��󫯾��èR�_|��-?�����'?�ɏ���^�G?������ā����wn���]�������r�Jw�5�Ī�\ ׂ��?��g۽<OH�z�	�Ժcǎ�ٳg�	&Ĝv.��~��8۶m3� ���θ�|�M7q�D��[��V��|���Oc2��_�{!�?�3f��v "HJ����6<�x���F�>��ߚ5k��Y�M�����'�4B� ��P*d�w�}�<xp���	���,/�F�P-�!Bh�o�>Ï~�#�L�!R[��x��)�.��w�Aj���k����Đ�/	��'�x��	A����g���{�1��R���0֑~�^�o�o#�������$�HF��4D� �,���@���&��C�$��
�c=#t�bB+H�yݺunŊ���� YI�>���2$�>뺞#}��߷qùh	�D<o��Dt!�z����?�uO��Z���On���ŧ��B1.��o��q���EN�P[q�@������[��dو��G���O2�W<�LG=K����o��O�2%�WD仟�����!��"��P�K�,�qqb$���{�u��\�qi1�W�AyL����y5<���!s�I /��r�!E	9���`!��*�/�T����� ��<S���,���*T�|����u@��D%.�M�I�;v�X7u�Ըo�[?�~u�� !p/��<y�khh�����Xi8�� �mĚ`z�����'$�:/-�r�µE�����tj�o�;}�HA���i<��PMh,���k�0!@ߚ��H=}���XT�;�e��g�R.��{�{|��RM�ޙpH�
yٚ�8��]����@�Z D��ZVaCD�/!g�{��b��Da�2e~2/�!b-޺O����f��<E±�����r���&�&+�^/�����q�th�i"R
�����j""H�j��b
M��U,!��Qqo�k�R��7A����%��@,cb����a��|�>>~�x�Pqv80:�J:B�8���{�X��+�S�B�ϡ�+����D�E�1H�>d�K&�z�bK�;b(p��IZd&�N��`�Yܦ8
�3�p����U�nBm��L"k1V?!����Ȝ�ӗ��z���ŢS�!q�����e=1�+4�����sC����L��E��3��|�N�pQ����7o�[�~}�0q��$$D��466��I��6�1MǏo2�2�C�q/�Ƹh#�S�q��	Zh�G/�z͂���ڬ���H	��~���G�����؈�sB�"�2|��ؑ,
u!���N�>}�ō'a�\*Ε����3g���y����7�l����7�"Ή'�1i	]�����5~���F}�]9"�v,���ImI�G�a��-���t!~��a��\D%����m����W�v��կ�4#��?���;�qn�O�.��N��>|8�0& ',�\�At /����pmеe˖Y4��	E=�~��&t,�G��R�a����@�BgR�2ao����ѓuv.b�Ջ�3`� w����5k���=e:W�����9M�h�$�'� ���n2u�}�����k�i�#MC����2Qi?d�w�}��as��n4ق
�@���ΝkQar2b��DE�}�;�q��a.F�J�jiҤI�%dΆ�袦�
5���K����Y�a�֭]�I8e֬Y��A������<�m����a��~�g755Y�ČP� L�
	f�0ɑ�;��]w�u�Y��0'���;�Ȍ���t}�R���ꪫ��C/�>(��:qg̘a�>*�9I�2w��b�i�5ɀ�Fy�
��=LN�P�_iX�+=��eR+��R�C_���4I��$�I����F�ZF�e�b.�*_C;Ƃ�����2w�x3`��7.^�Bs;��s�A?��$�-zN�P�6�����Dx T�8T\�a��"�0P�`�LVaO�Y?aH^bJ]�
̑�&|[6T�K:��������~d��4���3� �����(���Q��
-P�Vl!�Ο�r�B|�w��sX�z�g*Ǝ����SI.�T�?7Q�Ԓ�)���H�Ty��d�9��]���Ktͩ��OR�	#������!U��{����5����>�?���%�sz��:0�����%p�I%
�v\<$�i{��K
:׌�q?���L�{"��ޗ��x������@���ʟ��+�5�~W���*9�@�<�1��
�r��*{FY䀩�5��%U9�-�QyNo��%�,�Py�!�5J�<]w2PXE2DĳU����B
S��_uM��6�������b�R�+㠭9���mܒ#�rũ�Q(D��\�M� �*�u��!���QdI�#�����]M]��z�te)W���C ��4e�Qh'�
�r�2" Is�K<x0���3�>�*�U����P�T�L1*U�7���;��{I!�c�*���8_I���*���cO�oVxp!�Qۿ���(��p���$"��e; !x&�\Tq Ry�#I�J$�~���Zvr֜���gM�,�WiDVn�JD..ݷ���T��:or�/�0/�g�H�EWQZ��V�>!�J� D�ЎRSr$�@4����=%�2J1U��X>����LG��[��{ ��l>eDU���{��,�d(��%�ѨE幪씂�T����[׮]k�@<���x�^TR�G�B��ח,����[o�ĭ�}�e,I�E������2�!ÆZ�I���ܕ�������l�J&�vt�%���VKK�ۺ�uː�=�~�{��o�"�͵��ߙ3g�={���׌rC��~ ��6�8p��
"�qChCA����]}�p�b��8xPA�{/2T2� �m��%���-ɓ�e��п���4������!���K����-��3���\����z5����>t0���w�Ͽ��-�3ӵ��6�Lj���7�=���u�g�tٜ����Lr�{���~Teu��䲱��ɐ��Yo\�/�5E	&"�'#H�n"�إ�g<r�t���D)�L�ݸ?m�w��+w��Q7��1��;ݚv����)Mn���,���6�q���
�O�������A�P�7߲�	|�Q�ʏzʹ-����]qzę�m��"1�r� ��?nv�<����?u�7}���gǬM�7?Ӟ��<1޲*��c����F%���z���Zk�[�:0�EPu0&6����c�mϸ���#zw���7�|���	�QW��b-e܂�F9lOr�_~��YOK�9�._�J��pʪU�\�R�lڕyih�D! �N�����i��8w-��B�?R^�z
J����j/%9$��t�?#�Uo-lCO�旕E�u�_��"����J\*j*����2h����q�\T�RQ~۫��BuGڷGb,7�ѷ�.��Y�kkj��)�a�L�����k�a=%[��	K�YK�ٌ�'�d����{,���~�%Ӟv9/��^����W�L�>�/�I�֜�D�j��_�P�������	-ԅ���D��l{;J�N�<X8-.`����Gu�«���W׏���#�ͬ �n7�hoosuu�� a���Oƫ/+ K�l�roiy��F~MMu� �#����Z�p�
��(:�W9W	f)��j����p�@VE�IS[
�E�_Y+��f��'g:�	tD�hL�ϑϟ)���+���jcK"���"`%�>*���K}�1��nB2��zJ'AMS|c�C��"<Uf�����4r���
3�ۼ	Lm�ݓ��PQZ�KP;������ٔ�0�W(��(QN�2.�Wރ��!8�=%�M��!d͐���/���'��ouw��*� �p�so�����ȭ\���-��o�!��_$U~�n�kF"Q�i/�ӱ�� �����Ϩ ԓ,9�QW"� �ғ��L2��Kt���Hw��s�d�O1b�KU�Y�����qo]�J3o��Y�i*�Qmn��Jeɲ8r�.�~��d�}]݀x���wUk��!�PD�<�T�C�eO_���ү��}n�?�3��z�U�7��%�-�?�v��e���G>qM�]?o��kN��Q�����]Em_ˉ`U-�7��0�#��@md���.����Vݎt`UQ���X/t_OC�$���8�2��Q�2e:���xp����N���T�#���}����c��{w��w�r��Q\��sn�࡮q�w��c��j�Wko�dew�m���w�Y!+V��>�~�Ǉ�3	׭_o{*^x�E[��Λ�6l\�v��i[�{�y;��|ꩧLjz���\p���=�6NO%��9v��G�>w���.Q�����͜=۫��Q�M���@�J/1�!֏r#G\�9:j��nr���we�;;��y���N�~�@B�F�^DoaT�� �$z'f�PR���h�&��wB� ���6;ϢL�h�G�!�-�Ȳ!l"�.߽g�[�a���ϟ^�;:�}$@���3�j3�9��$���<�b�n���?��P"�HZޢ��d�TP[{��dN�#�?u�f�qS���z��5x}��ڗ�	���ܒ�f+���l���۱s�=v��9=gQ�T����zc����%n��]��O�'@�~��d!��<,(�P��m���I��L@^��B�{J&��iKx'���]A�ư��n�ĉq<誑�nrc����n@�:��kK�b�*��^X���\.S�n^���	oa2��q�/%Y���evϢ�o��������b��(/�q������TR���܍�n0�<��GnJ��nd�	(�5���6'fbg�x�G�6��WTT�u$ZoI��3g�=��O��&55����SWc:e5,���[�'����%-�qӘ}���Mf+R�G���h�&&kxTPX%�}��ᓪB��G2���r�-�\�,�<�%e!y�*��.a�	�	���\FuS�t!�W�W��%���[�3�=�L��μ�B�'�ϷFrՕ�r�j9m��g��U�O�V Q�o����(1,gQ��TD�ɸ�����Xq$�=iY4��E�,�$���l�P��,���;Ot�| {H"Ý��La�'�d���ʤE�-�	Yx��%�y��ݝ�p�T\.O��7��a'�������(H�鲱�62d
��ITHݫx) �v�RJ��w
�l������F�

R��i�o��g��րT2�;��w��C>	O�QWxBuXoK_�����kkF)v.1�� ���&|��Wv��J4-�1VeZd����;�w����V�iu��$�f)�H�[��M��Q
�ˁ��X
YO8}��x%��p����pb'�3@���3i�S�P��H������H��D⽪�oA���ٶ�J�N,�J�ړ�U�?��TS%���Ų:�[��#k+�IX���:ᐝ:u�͙3����Ǐ��ߛO�0�z����m�����z;(Iz��W��k�kI�����Ĥ(	՚E7<c�"�.��^
!��֖�-%28���G�#��M�a1u���{��C��'�]w�e�C(��q�3���d�X�r���w޵ҝ8�L�yw���/_a���O?i�%иs�N+�$2���/F(�5�)�]<�9���kGEEtJH"��i
��GP������������qc�����YQQ"��
ӈ�����F�⛞K�P25%gK���^��S�S�PU (*�tv��8�[>�� �8i���w�n;��괝,
�%c�AU��?�`��B�L�Wv%#�=��p9�BB�  ߑ���)f�W �55}��9h� �����)�cMOzuӛ�l��9Xc�6ؚA�j�����WZ�!�Y��(�d'$�L��ڿ! ��-
�	m�EmM�pm�GL8�Lf)GWs?�­[7���A��Q� [� 9�!��6�I��%[3d�k��{� ^B��ދ�ů,���V��%� �L4�n���g��g������剨�P*�������B֝���Ro@ɬ)��������:| +����!�N 0�I��rmV�H_XQ�'<K֓�g�	1�Q�{B0q/�d\�?:��.�#�.!�$FG�'>�@�A5�;��+` ?Oj��sG�� Q�㻒��3r��������)�n׽�֜N�M31�StJ�C��ct���_��g0�۶lْ�T��_�����,l��kF��+W�z��_�?ަx�(-t\�/��q|ڴi��iӦ%�J*��J����,_�� �bbx���_��ߏ9�`q���P�A�?��?���~f׺T�L�4��N�8qݩS���VY�_xf�dԨQ?�]��x���ڵk�v���777�}��+P
X�	�O���������r[s�$    IEND�B`�PK   ���X�\�]�� �� /   images/8e60f633-70d2-40b4-a331-b1224c91635f.png�y<�k�?<�(!uJd	��B�ĄJY"R�,��lc�c_*T�$dK�성�d+KٙKd��e&&��{���>����{^�^�ܧ��}���������0�AI��l+c>A�|�G���؜S�F~\��?oG*ް��8�A�PU�\�
>d���e{���u��.�B	� �ln#�
ZZGN��`aJ��^s����<����w7�ο?%E�����0<(����3T�laй��h�k?�]K�����!��n,:���ԫ�=/y�#�n��x�~�U7�,y�G��L�(�̛?�?�����΁+��4ٻ<���Usu����Ȇr�ӧZ�q�`�;�+���-�GGG7%�PE��݌���X�dK�W��	n�0����ƕ�I��"ia��q�v�����ТV��3�"l�-���K�t�@`,�>�鉮��>F��YeV����(�]������A��z�X�xx����w�+�}8�JC��\`s���<�Z�_x4|��|[�2om9�1\䶸0�+A-ρ��W2�E��̹͝��i`}�>��Ep�Ԝ���T�g'#�Bު��}6�\������ڗ��ʗt=-�ӑ��i�Y��=Șd��%�CXC]]]�UK�S���e�.A(��b*J�zrr�f��O-��v�����/��{�;��[uӺ&��9��Ħ�J��d������LU���酸��3����fv��^*8��շ	Z��m��z��@.���"��&˓���?����)��^l���"������񽬌��'~J,�����o��?�MKE\~8�KJ�#%j��$��Z+�����wb0����� ���0��2O���1j��i�з�0U�b���&λȀǨ�3�b֔o�Q==�3B�5{��Il�TA�p�ϱ��B��]gg�,�~���|���`}<��e�if������ľm��R�/.��6�\`s��6�\`s��6���?k8���9S��=勞�l^7������u�yݼn^��w�믳 ��ϲyݼn^7������u�yݼn^������?�>�Q���N���\�x��qIq�ș���!=8��;�%x�n��'���d�A��k��7�խ;����y�Rw��`O�p��\�d����b���|�ˑ���I���l�ƭ7o�Fwp�)`ԫ���6?��`��6?��`��6?��`���>�H��9$������uwk��>�����.�w��Ǽ]^�y뾴D��蓻�\��<Y�#�L����vn��SH��r�:� -(�����߻�#Z���e����h��J5�N�/���	%x��y3��GG?#��4���7�nsiƖ�7�be-��:�zv�`���E(��댏��e~���>Y�L�S�Ll�F�/a#l�����/+�'f<����-��$73<���r^>�K��-N�̔��w����@��6m2mF�>"õЂ
���{�Pt��@'��C��[�4�ǂ�y������2��!-M�W��]���F���ެM����:S�p7zxF��Uؾt�m#���e�佌Ŵ�nY�ö����Ȍ�^ӌŌ<	�[/����ݽ&�3�_Y	�?�����u����K9M�\dOYL���vҰ�y����I?y�m��8�����7��W�&�*̵�v-,-fI�e�ĜX����}]s�iɒ�j6~�C��6���a�a�a��5/��=]��z��=��t�4F.��XZ�)�C�<c)[�E�e.�u0�.V����,u��h��X��A�]��w';/'/Y.���i�ʅ掁 ٶU	u?��o��C�������c�E�e%9y�)t�I:�a�S7;l�3NI7N;F�5X9FX�M��V��������\��{�g��<��.�.w��O���нˋ�n�{���K���%�..�i����u�H�����Uǲ��RSYK��J!N]E�m�BA�GY��jʹXњ�r��:�5�|���p��n� x"����)�P�2ۈ������T�*�d��{��
��\���7�t�_�n��ji�_���Х2}p�[��c������3�q�+�Gm3�t�
S�P�1w-e~&�W3���y�h�v�U��)9�8�@�ϯbQ4����ru���F��a���Mi氖^��W�99OL�(��V�*������17��n��)��R+��u<�g�p�1��"c�D��Tno��zM�`?-�~mS�)���Z&-�2��>td�[�vp��zK�H̽������ ɜ���;�K��1��j��LGk���&�C_ƣR�M�����J�F�]:�}Z;��An��ȴۈ��,���v���Y�P�r�Lm9?wu���}x��I�\�b����v]�E�N��l�!�2f���f�[�w쥰Ms-��S!�3,����㖣�����02�y�
��G�<�ᙣÌ*q|�S`�l�W�!�%���T��lB���+,�Ӷ��!�u_��]��������"E*��8��͢��3\��ID�Y�ϋ���L���ˡ����K��&�^�ʗ!أ[K���;��$�;]���-�zh_�,G����/���`,=��U,gMÅ�;Q�~�!�l�=,EE���)�˛#ɐG;�rp����HOr���2}/�X�?��uB������A,�]RI�E�����MN�����"�S��8{�"]g�p!\��'�P{�i��b�"�!���Q�������SB���;(��2��n>T�"� |��1�O��G�|vAjm��G]ـ��(�����&��Wx�uʷ�:�ZWd�Y��j6Ё߻���e������'d�a�����2�����)�g�2F��Ua�~�0�-��������!ݮýE	Y�E���W�٪����Q%
u'x���c�`��ͧ��Bq.=j'�e���?���U0�wd���!X�*����-9F��^��]v4�:�l#d]�a�"��R+�
.������C�25����h����'���T��-��`߅�Q���C�H����������T�Ƕ�Ĵ�=�ó�u�B7��5���z���%wr��W��A?�*ݮc��CjvV3��"�R��%<_�!"[к����;��R3���� R�s�֛^�|�Q�s^��O�
�&6���@;���d���c_�5����K�v��-�7t���ә��1�q=jD�pWr�ntK[�����G�h�z�K"Om0���t}U���Q}�ɯi^w9]����:�}���zfj"/����S���a~mR1�\!�>�g'�Q�|�W��o�z�Op4n�3�ݍ2
ݚ�~9i�g�)_��������
��>+jT�T�cf����B��m�i�����!�h[�jb��ѕ�u> 9�=0�����$"�ؿ+��U�y�x����︐�~w�x�V5uޕRޥ��+h쟜�m�ePkEM����s�"\d^��Р�
y�G��騰qƖ��\�a�K���pj�KvPHJ(������Ř�/gR�*���|d��r�P:�畵	�MoU���`eF������E#�j���H�{ej5:�	נ�e�%�jouʦ4��b�w��`�]$3�yx�O����+���~���'��P?�֑�(xP��$l�YKb�Q�NԨ��vJ���6}�����a��G�%��~�H�F����ė�mo��>��d晸��y&mU�����yM7��w�����E�6h;p��q�D\	��r����8|�oE�Ө]��_߫��#>^�ʫ���-b̞�U���!�DX�������?}�ȯ �Ǧ��/{�¬w��/�5n���Y���������#f��t'w�[
,*c�p6�r�Q�ڧ��w�����';��������B�g�����2A!��SA�Bu�*+P����������[�,�	Yŝu0����R��70��F�V�ӟ�b����	����NT�>,�C���"WD��_Ң�u���%�ip�gѿ��:�)�zg@C��P� :z%���/ 95�=��I�����p�G�1u����į�e���H���h��/�!�{+��A6x������6����y��=�{�KA-�ß�����R%�5�x;]�jCFj�)Eي��3���'s���)6Z�~�5>�i��>k6��6���iO)B·���m?˙u�5�_ɠ�����%���2�]��t��"ߍܦ�<���?pb�ó�+��1����[�A-iB� �R��0-��Q�T�|�e�k^��
W�}����Ϻ����Hj���I2�������t���K�e�
©D��J�BӁ���`P1��c>�	���Ev��$1���T�.�@�ȇ��u��oO(����x	v�X�r_9��@��d���ϙ�H8����c�plŅ�~,#U�����CS]�.B�oY.������ut�c���.��gF�QP8,�"���e�I�bD�#�D��l������-�[�;��y�[�c��վ����l����PG�I��D�	21C��q��\�!, ��2�ң�+�>~C����X�>��m�*�n>{q�h;!a����&���Ə4�HT�|vQ~̈��� ��?��ի4�"i�mV�{)��=�$zo��4j���k���'cX�+����Y�6۱!9G	_N9Q����b��xN�v%��+��vO�g�`	%)�ݫ2O����Ե45ik����u�U+�ނ��%ykД>��@��%�1��a�E9&j�掎B(�ӽK #! #��Ƿ\kk c�[�� -S��T��B��"D_���q�^	�Ğd>���o>+� �Xy̥sPC���%���ȇ����^�.,
}1�����Eb	��э�%���Η��@H
d�0E����Os����<|��)V�'����v��}:k�&���|5�Y�Fb�'��Jg�s+�� {�b'�������}`�J���+�%|�r��G�%�-��,I�	G���>��e��[Pa�B�
5���;#2�H3�9���J(����x���4u4bn?�`����7(��kK�.�h���5$����U������W?�[�����o�j�*�++�Y32-�[��?�/茱�*[�V����k��g@{�Ԕz��`'��8@����
�L��A��kB�eR�
�n!�m�c�'�/r�ԋ>�I��>�9����Hwg����5r�cv�i]��]h�=����0+�GU�Cm@��?D�?R�;���ŚϸrN~8�>iiP�g����Ѫ��+�����6�e�4�r2CD��ԄĽ$I�+�'\3��>�be@c��Zս:�/zCX!tQ/p�J{z��D�S�a��{r�SğB�)K��na�"y��!O�����Z�F���H�F������bn�@Re�Uk�.��f�Gj�8�`��_p�V��-���,�ó�}�
H "����M��X�[�^�쾊��mT��z�y7�����f��:�3�B���2 �����r���q��0[��4��?Q�[;�n��mtX_��D��9j�g�N~Li#9��}�mף~����S�$�y@z��ޑw�o:a�s��`'o�:�fY���x���f���o>+m�xe&�Pȏ��_�n��O���F��n��@���רđ/�Ɵ��
}7=�_���l̜"=6�6[=�r���("�C ��;��_��Z_��W"�X�u�:Y�b$5�"���Q�*����%��tQ${$A�\����A���y����>ƒ�70��v��O@�� 0x(v>[f� �U�ۗ��/徘Vs�Is��/��E�˷�����g�<\a�Վ2��g���s$�7���m���0�?�,*��I �]�"�֌��S�S���uٛ�n�K�(�U��wF+���������9��p�_k����[�#Q�b!ct?�R�"F �qE�zȀ�*�aokܼ�$Z��F��KI��W�jv���'z�a}q�o?xmڔ�'3�&����5l����+8b.�.y�gI'���Tw�PI�����<�4������L
��x-uu.@�4�]6q%e�#��0���Ӏ{�`�����1Oxjćҏ[wQ<+d�>C��sP=K��*���\Zo�D�!�������?"�Dϕ��@ppq�O���Z��������C�U]��P��t7��� |���T�vm�씟��:0=5��z�|mu)tln�T��%����-�]�D*�o*���2a�NN	�^�ӌG������a��O����q� �h��6,�ue�0O�zT�آ=5�ǲ�����^�`>�E���E��p��T��
^ɵX+})ů�%������@�.��G�Oq�65�޾�_��vتgm����:F�o�[�F�Uj�o��s]1�P��c�e��'���[��fk뇎�~��Զ��X�;�ڑP�=�U�k�mt#z,nQ��j�{�o�� �%�(�ͩ(�T�e�k�tr�ܝ�tآ��|!;|-�,��J��9-ˌ~�)����s�r}2�����06a��l^�(��V�Ę�4� �2gx&����y�L�xg��AA��3K�R8�	��S�K�H+�&	4W@un����Z��A�Ǔ�W�:k|��V�Ʊ+e�F=�:H7[l�Ƶ�L:Ws� ��q��*M%4D,cg�Vp�h�/�o��T�k�\k@�(���
j!�7c*.��|V&*_]�("W�G�{���
�`���O&�?O��P�񄷤e��}(�x7o��pxziM^mN�kVDs��&\CG�(�����po�"��t(�[ޕa��k;6�[�J �\�f���""$ț��ǥ~ž���ɉ��>�w�9�łź�[��w`j��h�/̉T���x�v���X�-�ğ�A[t�6��Q!L�f���=^S1�4@Cp9�)�C���pM�W��tM�9���:��M�x|i���-��E�Q�׾]H5�u��Ĕ��g|�H2 !��55�|G]�}�(���~�uA���8 ��a���Ƥ�v�߅�OW��-K�R�����h;�-^]w(�+	��������]�_K3�L7��c����+6w��a����g��hOT�\񬐎S��i�ܘ�+�{�젫�bBb�PǏ�9�<3���:�i㵚�@ھW2�C�co\$n52GU�(�kjw�����iN�����Pb��'�#c���o�`�Bg�%(3ªǦ_]�@�7_�r��c<�o�O��~N FT?�I=,r%l��s�/k �����L,��f�gF��%�$�EWYx�'��q]������Y�^K� �11�Wꖦ�G݊���ƃRN�S���B钤��j�,��E��	 [�!�M�1�U�x�Ϝd�x�Z���Tc���>�k��f\��a�F}�0���4��:C	%�tcc��^�:а�n�Q�+��9�������Ξ�F�k�ڬ�S�Go	 4�y���������./=�E���A���z�[A��}B)�KvzUS��T'�-X= 
أet����W�+��>|�E�ߗ��젴!OÇ��N�]���z���K�����ذoNͥ����מ+�]�
Ch.�p�G���4|��Pf�����3:l�?�Jǣou��c�)��}
+��1i	O�N�;��q���]tBh��m����閂z�>�u������v��X�GFR���<2��r�^Տ�D8c �=^;�t�|��7��3'�f�����{�2�� 5jD��?�j��1��pS�R���e���H�K����Ж�f�[gƆ�}/�f]�S5ٻ/�3r!V�50*q���Y5����4��u��7ƕp�$w"��C�Q;�4�B˺܆���Ԥ�ot_τ����Z��{�+ �SԨL�%��r-�u�cl��\�=����'�C������b^ɛ�aXx�$6�դ��:s�_�O��!�e�}X�[;J'tc#�z�Dde��kM�Z\�QtC]`wi�BE[�����8CY�|ן]��fk��12u���W��4 �g#�W��>�B�	kH��叛���0���Vhj��c$�̏��<���+�)թ�u�\�F�E��vdE�U��|>�lh�xPT�v�9Kb��k�C�4���tT�sf��	e�{���Cb��C�ֈ�rﶬ�V~.f4K���|�q�7�׌����x�@ְڕ�B_�	��+nD�=���>/tM*ɑ�-�?�����N�z�arE�[	�,�X���_��W�c|<J�
�������"�1���3�g��UH�:���Z��c��7��Fy[�5<��B��]Yqn�}��2�����}/"���A��p���� `��>�
�5��b�		����3��^�J5��?X��@�l�n��9���tA��[(Y1{�\ӳH�o6'��q5�����Xn�ա :}�@���m���쑤��p��u�J�IR�P�l\|�M;-SY*�i�&߬XS�����=�ƕ��&�S�pM�{��ޜJ��+4C�Ĩ=O��L��yB���Z�6$'h�5�,(�F�x�b����9c"mɜ�o��.j�Л	y{ã.߭|�0�7
<���E3�<@�{��J�)����5D�6�9H���J���Fn{��zI沈שDXz;^"
Y�3�W�9v���62��+\��F��"�����$Ϳ����% Q0! =����㒎wU,�P�n�4���8�ƀzn�{�NA��i�!��E-s�S�R���	5��;I��Nq�aooAx���"�W�L����$,��W�+z�����GI�l��w�:�s]Lܝ^~,�i�)/���
mBgq!��5���?��J|1��_8���>PK�����9��k���}ݦb�o�F@��~�Pԗ�b˔
�(q���5Qj/>d��kA&?�@O]�XL��9E��In�b酛Y:���&hчBo��AW�B:�t��i���ZqtZ�d��ñ��91,���Nt�\{���V9f�v� (}�i�L^�#FW�K���gQ*����`Y"ߨ��e��k���5+���mB�N�B"���5N3��s-�i�|l{�p�@W�����\q4����>���!��-��qX W���!{�/T�����K^U�L��<X9��,@����V��'G�R�j���a6BB���Y~V�	+�e�L��)�*��c�����6.���Yn2��V���
)#Z?��B�!q��g��/R��L�r��ڐ��M��4:k�����4�(�tz��K;�K8a�|D�JZ���282=��q.i6�D0�:�9�~*��33�R,��ʒ��]i��D��8���_\����(�)�J����IJ-�;>��
�g�mFZ�`.��72��]ҕiQjY=ޖ�gꏁ��%�%`H'��������'}|0���y�i9����5�S@�ߋ��X�P!_I*�k��N�gT
��0L2�?}׸Q�8�5��4���e[awΗ^���s�{�E��|A4����%��Ep�c"Z&#ɃS=dw"��)�+]�0����;���/���8���0:���\q��Q"&c(*UD�Z�J"&����ړ�y��X��.I�����0}O�0�w�:�� ��8[�X0�3-������ϐ��u([��%Mi&�V�H�k��ԩdҺ�������)s�H�p���b�l&h��$�X[x���.���U�b�u/����!%.=;��cM�,񏜭�.����YB+����%��n���M�8[Or�Ur�@r<ͷ�v?�'�y�˻-)���pnG��?���H���׹�Bwf�:�r5�٧�YW�4����FWJfb�:�(Xd���?��`"��=:�.	��Z�@y1t�{u�6Q}?=w��2嚨,|dn}�Ќ���Bjp�?e: �@��}��
 u��bu5L��?��S����o*��9l_҆�M�vqV�H����>,��4#��Xn�~��k�q�qŮL��3�e�/�LЕ���zʤ˸U�bm?]����[�扱�2j����r��.<R)��	���ߣ��eCG �}aj����دe�)�2�k�|�_�H|��Ѩ��+p�L�^��_Ɣ�V�f�>����@H�e����� =�A4�E����a�%��&�3�i(}���g>�ĞO��!�O_�
TE�ɖ�n�Hp'&�7^����ˁ�:��A�8�nGC�n�%.��`�����j@�V��!�$pV.�y�/o{��C�7������_]1�{��w��w����ߺ�:���y���� �(�;��~w-ʌ\*��<�}�u����^I[8�_�u�f�;{|=Ń��j�>�&�ot��#�W*l=�xP�	���;���f�Ptw�(A,�c�@$g��#&=�7��VnD�ƒ|TH=C"!�p�p�`+n��V�Z�[��d9�v"���)P�]��/H5]Ñڪ���O3|P	,y�R���v�Vî����c̦{��.2���I��T����U���'~4v,x�1�>�M���������D��N�	6;]�޽�<�@f(1u��}x�XhL�We�@�tk�oV�e{kU+9^�-q����z�9J��sA� oHg��Ő2nJ	�^�E>&M�%��f䰅`EP�/�h�w(��f즏��X
ޟ}aW��-sw�7<ծ�^�c{%-�����b�t����_CČ�����1���B���",�R�[*T�_ ���!���
S#�٘��NH��N���;⋃�>W�
Uw3Vԥ@��SV�o�N�i���#�Q`�hp�=�)P����Q���Q�"��<{�������js�ЎX6xR?�g_���q��:=�0��C�i��������;��@�O�(�x�3�B�\>�u��H�,��7^��z��F�£M���N<Y��s�$B�y�ϱ���Ƽjhѓ�,9��t�����@�a��qOE眾�7��1Sd*��H[g �L$Y�8 #]��E7&!`�yX�B�d7�;�PA�j��V�������0
l$J?Z~'zZ*32 �oQ�}��]��UGx�|l��¯R��9�[�.�0�����z�S;��R�6�خӛ�Co9���m��cl��:�xZ�QoP��VF����)bx/(H�}�����Z�V0;; �� ��w��<�e9��-'��2�s�s���_�`�C�]�'aR�Q����ܛU4Bk�n���8(�F�p�fԱS7��@S\�Ѻ0~�l�A���c}c ~ĵrN{��j�o_O�������V�yhP�7��1"){}����{)"t�`�V���c���D�Q����JK��7F+|����e��=�^�C�z��~�n��	JQ�5�_�E@���E�@p��������ZH�z	�aMnW_���S�������`@Q. s	�w( ���͌���A��J�*�M�|�-�5���Z��z& /�#�|�	�����L�/�«vtٖ;@N��D�7���C �N	t���E>�� x9�*��a#��[�i`@�!Ѣc��������JVGI��-H����Q�v�{�ڔm��7���)F<����󳽵���g�v���p����<� ����}RxK�a�U��A��ߏ��v�2�����D3e%���%�"���ޢ��W:��^i�T����	'׶W]�ޔK��[�+馤VH�2����U-��BP�W1+�x3O0�ka�S;�R���8>*J���տ�!S��u��_0�)����'��nZ��,+h�[٢-����v�z,v{L�� ��ZM�Llب�i��ʵU���	d��=�M����}��x�����ǵJ;��V�C#�ܒbX���[�m�^_����dS���Aa0�pB���p<�y`�nQ���"'���������%>G��7r�9O�&�sk���O(��K�R�]yԽ!���`#�+ߏQ_/cU.lφ���EkR����#��!���7��G�Ǟh!�E��K��prI�Q&�%���g�K�.IH��{mMw�0�������������&�����~1!���`�Xj*	J"���
/��L̼b���wj���2���7°�L�h�Ⱥ����ojW�I�����pn�c��Q;�
V6 �o�?/�o��L�ӂ��	Z�S�u���c#��&��uRt5���*~e]��Y�U5��b �����	\|��-�<�/�鍯笘0f3-���`m�<H:H)��T@z�a�.G���	2@����.M�h�D��h\�Y���] 4�lK���s5?4�S��6��x��	F����(�z������ݖ��ZUK->�p�ҋ��t���Ї�h�HG�3FW�a'� �<��??�MO,d��ݜ�+W�� %̇+'�
;6�Uj��AP}׺ �@��y7N֣a��V�mr�e�\��ʿcu���ƚ�"���*�}��AF���P'�o<6��/O?���@�:����:�U��8�x�ϧ����#=Q�!��N>�{�C8��}�^�3Q�#Ҿ��]q���+�[H�ix���@=�3�l+�Vz������f��t�<��v��������\�"ȍ�%E΀�Td#���_�r�������T+g	�qP�K������H}q;J��2����*���V�5���]~0�|ݸ�V��Xt�j�_N�C1��L��28� ��F��q���t͉��Uq���>�����L�9�qx���Y��d�x�0<J��v��s�	p���rV��T|爄�����5~��������K�r�����������\f� ��Bw*��Y�*]��|G=i�cx�|o���G�<������#e#����W#�߼�m�"�t�Ħ����w�8C�xg���f$�)Pѥ�3"��\����1�~�>w����p]e��TL`@��&x�Xt-�dt���=��$����{h��ߨ�nOkH^�����{�o���j�,����Ӟ�z���
�|�z+�$_��Ȱ���JD�P��Tm�����Ǵx�S��	��mq�=�C��x?3jD�+�Qu��$M�i���3 ��;�E��K,w��Y�����٭��w�\�Ć!��G#�w��H|��S��ŵ^[���^)��ޛ#�aۧ}���|�@%���_��#�uT
�U	kz�e,r%��T�*ٯ*p1.��y��{�����$��������j�gŰ��`'�g#�̙O�g�?��4�=B��F�b4� ���w8 =��Lΐ>-�� MY
ǔi���]Cs1��\qV�\���b/кU�,�a&��޲����Aѥ� ��d=��옑87�����
�&��(�3�w�rş�ϝ��g �ׅ5���p�FL�LaH��Du���~=�Vӽ#5�)��������{����ϰښ��[�sؤ{E�s�)��g��D�{�u[��s<��e^y$�gŴ@��2�g�bD�l4����I8���祷��}��&h��oԟ��d�l�����.�?U���y3�F�>W��|т%�ëc�t��'�a�ΧPn��6q��A9C����L@���H$�@W�T���N��^t�ϰr�-��zԧ!�R�X:L�����9���(�J�+V{���MG?5^N;#%V�zwӇ���G�9���E����l-H�[_iR>�ĭ'�S�Q��,ü=)�e�G�9jU֏b^��֨�hU�y0n=WM9�~����o�PU)��+X����eH@��h=ۮ0{}6�C�k����#H�=y��{���ж��Z*W�F�>�u�'Dd�۴���J7vKï����x�мfԂL~�*qQ<��R!z���[�R��x�X���g^씡n�5��H��J3�n�?W0�� �*5�����pYm�7(�14N~��OU��^A��X�SUe������>eP��fQ���'�`@�jB�����n5��4FFj�5Q�ݵ�p�("=1��ɒ�1 tbz3���W>�:|l�_{�ߨc�=�e��p�"@#� '�"�������xe��OU�)��Ŋ"B@ý�i���v���bXOۍ���>��&�:@3��p������k̷��_tW�b�ZqY�
��ԳK+y����`=E�"���t���D���d@]��2H��ym򰈱��5�&V�;:�̦ ȯ��C�ʄ�f�2��O}�����C�^�Y[��A՚��U�iO�c��	�c� Pv� ���mj�Ϟ�?l��D�/\5
 �g�pY+.�}�����ࠖA������1�Q`�P]
���@P�8� X;E���|ihG�7�q�:�����"�%�x�K���D�9?����u�DS� p��=Am���G���|���HSW�L�w�:S�Z��U�x~�k�G�)@�a�蠮l���I�`��uF������62;'jX��_y�h�h�f�.Pn� z���'���d8/�*l��5OZ��֏*�������wy���^���ztP�uZ��CK�0����'M�&���f�-WAW��D�!m���`�Q{Ng�~w�L"�����S��ۤ�����8�o���5���6����-I�uk��{�bF+i;�ތL�t��)��s�	����C{���g��ݖ����WXO2}UZ�a%wڰ�9�`9��'��e����ԯ�A�6b
�Q��H�7����i�)	��.ΝM��H�$RI#�*��[��-�Ю��JE#6����΢Z��,[�a�\��)�@� �!O�p������a��B�ˤq����zS�2�$��m�s��S��ʿد�Fxc �.�G����"&>Mhz�q)�Ǚ��ȣ�a���|�W� oxF��1dM�o��Vi�[����a��X(��>��ϱ��y��@����=�����
���F��/#���D]P8<�ʮ��ʖH)u&c���G�/�M��x�]D�����Q��BJ>��y����u�ھ���ƿ�4�`���hy	 ���ך��|d�������J�W#��v���o����ױE;�Ԝ�7j6��'6�3 ��2|��;��]*֕��خ��IQ��p���x�$���k�:���b �
݅g�LЖ���@��j�#�U� u���m�,�d���W�?3PSW=�����:�r���;��Ӊ)��M�@��A&��ÁH��RȚ��?��aQ�����|�D��1G���li���������7oM�Y�z�((P�+ی߾�fI����Y�����P�WF�~�B�N˥R&K6	L��S�s�C���3�^��,m�jj�Q����>�_�Nv�þ�4�5�~���)c�Ŝ���@�L"~ �x��p�gTl!�O���ɶ ���Y��8�Y횎�8�dnDz���wIo<|J��55P+�B$|�w���Wz`�-���Di鴛A���`C�M��Ear�snt�	�H�|�_a�)�f�4됆��p�j(�w���BWT��
�Au��p"����,��iP�&
���l��֙z=�Vup�Mee�JG6B�yuU�V�Sw�CYٻu��!�e��d���g����*�nr�#@�)������uE�����
�
�լ�L�̨��!P�7���* ͕,ŀR/>;?2�����n$�s"с]695�����P}w�/*��
+%�����I���a�~D�.������o1ʸU�y��J?+*�Z�I�xD�R�l������KA��-sK��@|��5A4��[�JdLC��j,s�Нp�����u�ަ���Ͻ��1�o<�<4�)e�Y�F�Bڙ�pɝ�p�$M��-��jc/h��)��dn[��� ��z3ҧ꺥"@�g�F%����
m��Ϟ��$�t4��v>�'!44��xD)D"$��`����=o>����Y��	I7[�B�	�.^I��BX'��ˀ�4�u�2��%�Y���Ռ�%�8d*Y�O�g0w��L�ԭ,Vz���U<W3��q+i|�"����-�5�Kp/e ���9��@yo�:7
��nC���M�3D����r܂[&3������/|�Xd߲$�:�_�[�����8�v-6�J��)փ�_C��p	�_}[��sᨨ��Sf���i���6Hf)v>��=�~c��$WL����%A���&3�QY�+%���}D�$%b�o��{;߁� ���Qd"3���W'�u�8�8a`����������L�4��Q3�lb�T{?*�i�Ň^``��D}��I�`ilr?c�X�G��?���E��Nh�>�݌����O�p4\d#|_�^b��D��`H5y�_�|^(6��OY$��a�����q1lH]v�(4E�[����b?�V4��5Y6B�U������in�n��W�������_�<��ZX�Yo.ء�6@Yӥ�^Mb�y�ZY���H���V�r<�3�4��;6�+�v�H�ɵ�G�P�]<4�B������c�6v��_󷧣.�/�Y�����@o��QGC��}q����L�Z�*�-Y,�b@�;�n��FM�
*��L�L&�#�=$LЕ���(�czN�FM�s^¥�kd�j�(��0�Aqu�Ҹn�u���,�9qڿH+&�U�k�A�^{㿧3��Z�W�J��������|w�Ί6s
�˚�ݜ���$#��pݠ4w��d��P�L%�)��|����8���H��ߏ~���{�İqG)Y��k��)�u��.d�2��W���!:���3z�3����ñ��u�����O_^�s�!?�oX�Y���������{��q���q��}J�r�l��Wm	�
:�z�c0o�-�qEBs�n�|"8B;�Aԏ��h-��qSZ`(�!a��ݯM�7�@�u�t?N�/�No��V3]_E�Ȏ�l�Ig��F�SvC(�$���T˷�J�"-o%{�x���\v��_kuM~����"�Uz74m�D��:^�H�gR���F�|�!r�iC���׵�m�)�Y&h�=�}q�����|�u�M�ç����%�9h�K��>]��{�g0��a*ü-��5���!�m���Z�O�Wl��nV,�q���%��^Ob�ɳaz��Az�Wd�ni����i�k��`h���<��݋��P|�a$�,����M8[*�Q�����o�V"v2�ؿ�".T}N�8�h�1�/G�T�̐��OH�Hݒ�w��Ǟx���X����d�^��]K��s~A��t]�
.��Y�\+Ӵ1�]��/�?���g����6� ��
���z~�Pү��O�Ƥ��H��=����!�-^�0O�����s ����c�@��H���f�BB���+�k#2�0	B@�g\�;�v,�{��=�-3?�Mջ��[|�%j�<�Z�z��V��tM"dB�4��ho�kޤD�i�eY`��O�g{!����K��# ����('�:k���C��]w2�
4o?(Q�<��U/3X��F�+��"$�V�U;xy;_ݗ�@�Kr�{`꟝�����o?���ۯ[2������B��ҡ5��X/#�:ٻ�uSl��t�J��a. K����o�Cg��7�q]|��*9�=*�E@��=��G�^�H�Ju�	��zv����Id,�F1�t�Թ�=�@�j��x�|V�h$�E/��ܫ���O��g���.�I������Yu8�5�YK�E��F��c�q?=�@)����B�~)��Oo%n������0����/�NK��86ڗ䴟4�7[�]�IK>���,��U�&-�s��?���zX�c.V0�"��m+�9������?Ӗm�����TjZ�*�/���3�n������8�׸�&v���&CN��R��O�B�����:��:������X(Ƿ<f��Gt_�ƕS}��P�s�S!f�G�2rN�`�k�k�?�Y���T�勎���.��.�
��Z�/�C�fԖ�2Y�ϼ]|�i�=:���E5�����<M`�G�J�.z�։M$i.p9�݁"[�c;l��2,��Tn�������|��oXZ.��.Ƿ��'�4�<��7bd�Z�ǈ,�s(�e�Jw������ߗ�����2���t�x~n"�5�.�d�PH�ۅqY�b����kR;r��j���y���.��/��KoK��'����g�{��z��1������zI([����u�6�2���Qo.�{b�G��˽��dc�9&�����9��<��O�3������Ħ����ۥb�����a������N{J�$���F)�N��Th� K�l#C�崠,3!e�aD�a�R� L�,cHS&ːd,c���t��|�������1>�y_���|]�[q�t=��H������5������ͺ����q{�F�������
?�V �sO�<v" Ca�O�����Cs�zf�{�f+��+$fi�s#T�+�h�v�#h_�#ub���	퉎�w�kt��R����RE�縰�o�+BFP�Ũ��x��9�.�A�w�OصS�%��F����a�PHnd�}������	����z��*��DFth���/�G�$� 3�:�Vk�fb��d��
m.+y�c|��d��̈��(ڃ���:��9����ԧtwT ��;�� �W�ɘ�"��L�U�����T�3��O�&�.�'��	�??Ĝ��(6\�]�����ub�~U��T�Jt���A�ֹ��*#�m
i��h��o
2�(ёus����;�p�\��8�LFe������[.��W9�Ė�;���&�N�*^Fm�5s��Sfdm���V�žVQu�
4���y���KI��R�j� 6T�at|TjЕӳ&1�
yvH���9Q%�������Z%�/��X�ζ�W�f��j�G1ΓR*0x��I	2��(�"y�E2�$I���!>~����r��\C�R׎~���;�k����~F	������P	� 3��G��)��j���� �6F^v���fL���?$�/�%xr�
�64�m.�LC����jh�&�D������ᣎ��i�gjMXB�:|���5V.�4��Uܧ�ރhI�C������I��|1�k��fl��A�S���it�����Ol���RW�~��U5��g;i
ֆY�O�zm���!=�"d�sz�и�5���F��>J����gT?�*_	�oBP��ybW� �V��A��*��T�X������DI���U�'�^砱M�	�B>?-aRjT3����T׹��h:�ک�&tRQ��݀�x���co�N�GB�u���v\�湌��*���-�Gm��~���'#�+�Z:s��mә>��:���vy.7�
��0D��r����}jV�}cD��e�">{r� <[��
E��V!K[v۝�*+���[������o�:������}����	��h��������Hj¬��E��6�u��P�賍�b�U���7xt����9�2���T:����ٜ�tғ���	��t���F�9�/��c�|�7�}�4��-; �%�A��=�'��d4�ެ)��T,�.%��II��'�(:���UvmD��?ފux��}���P=�vyc��JG�CS��I悂�o�o���rxF(�7"��7
������0?ؙ!�(˴3��5�j��G��Y�q�S��|q$��o��<��>��X����6W�b��� ĚR{m�����T=�Y���5�)��G��^Y�>G��ׯ&�|��$�p��[Qj������ρ��hU�����w��w����|\��7\O�a�����l-?!�^.ȶ�#�����9b���|&��W��.�^�G$�
���?�׸�)�9��	F�ۃ�VI9dU��(�T�rʼvͿoR0��kĵZg�yV���B�K2�Ɗ��nq����$:��.���#j�QH*����VvV&�]X�G?����y�e�8�vY?0<�RT�h���9w%�X��ؖ�����_���A��qEKVk�!긣Vj�_馶��g����Vo?�y���Z�����[N?�V2��I��_�������c�>Z�Hp�L�v���/��]]��ǛF���p(j3R����=O�9C˝���]�9�}k�9�.�4�'�j���f���䙹X�Y^G:�mܶz�%T��t��{�v~}UP"5���+��DC�!:�?��8~�4y�KM�S皻������LGS�e�w��W�����nL��:C�y�����ʾ��Ŋ<���1#2�u�Vt�����Byſ�SE�T�"�}��O�7�?��n�9�J��"<��}�=	���O-=AF���B��R�m�FZ~�Ip"M%�D�0��Ә��J��& m�dP�ez�R�4|��"	#�F�sB� <4��l�E��u�p_�l?�̖�$��T|H@M�:X{�l�Bt_=4�e�q�T�P����F$�U!L:6Ϻo�䌧#6^�a�]�6h�|𡞩�4�4�d����9�mk�L[����<AB�EzHŸ ��e��[��jF$�=�w$p���H���m¬g �&H2�OQL��2��!�Nt=���=����lo��O+�.1X�J'G�ے>M��u|�8r&V���39z�pTL�v]+O4��Q��h+���_2�l�و��x]��>��c��p�x��m
���Y�@+�}t�bRn��D�v���{�RS�1}"J�Ar�ף�ӎ���)�z�h��^������;����w��8WV�Q]�3z�ybT�&X��#8Gi�=[�Q4h A]�C�K��[T���'e4`7H��<��� %��
Ҿ�:�1B�!�5����~�R��%Oe�:¶ȁ˹�D~��g�8:�k�Ud��W�ƴ����k2�"� 3&���oL��q�ē9e��1-A[�hg���a���G��ڮ�tK�D��w�-��.�?��(s��u�ӞV3ז6m��~Ǳ)��N(�Q�L9���ّ���*�ٵ;�$Y�I��#������� m�猂6dk�[�� ���&�󛒵�|��Yk�I�UhCO���P�_ ���4+���hO��D��©��ꎚm�8���N��<�Ŵ�3�Ė�#�]a��wz�$���d��Ҷ��Ì��P�݌�^�����Ù�sQ~�fv\��E;U�9��h+ �CT�|�do��'������W���DO��<��+E�e��θ��}iWД���Ou���J�q`�z�p��M3[�_ƫ/�0Օ���E���	P��T�Q������yq�&�ko�Λ��F��!�xr�[�4AA�N	�r������L@�̫r+�yp*q�<k���3"���M�b��_�T����$�+��5�5�&����#s��t �y6�3S�P[)�a��ql���#Y���y�|yjo�.���{/� Cǈ�ɭ�hR�
�y�����9���2}��X뻲���Ν�CΌc���m21�JJ��W<�7��.b%M�J��R��;��$�O��L��w3��_Mv(49m����躛��`,՛�d?�;��y;���Ř;B�ey�&��~w�|-��F��`�!�!w���	n�W���R͌�M���Z��k�s�2+󕃑8���L�ޔ��s�^���bY��:��P#�@=��~5���aH�k_J�������rXV4 ���r�H�X�S+h�6"i��%�l���<�Ц��oRKJ�ݻq�.��ix=\,������Ě�x�t/��U���c��J�	C@ ��sQ��P���Z{�J9(Q����$O�Sa;~��z�5~C<�ik��n`: ;��T���-J�����;t���Cм��M���������8�?�l��%�0T�����Po�,�J�VS���]�XvT+�5S�wxO�z~o���g�5?S��G��)�':�c�� C�4��lƗ�4z���>yvFM����}Ԅ�����<�}���G׮Q�'�O�$ ۘLYí�?��S�U������lu����|%lF�>i��"��eo����������w"���q���Z��e4[���>�&w�vQ�[�>�ki��[ך>qٻ=@p����@�R��X%(^[����l?g��r\UJ�	���:\U��'t�笉��D㱻A����x����K������.]��A������0�񠞲��~A���Ȱ��5&�7�y��{�̮C���ϖ05��;�&ib��s���(���SwRJ�ٟ����2ێ��5��Ą(�N@�r�[_sA6l��B�gs>��K�!4��|����Z`��GN������^�ȟ�f1\��j1ݲ���a����-^2gOaf�^��F��UQ�Z �q\V�Ce�p�����Fm�p��l�>�F�� ?��MEn�Rۦ�.t��K���v0{�Ka�9k:��bW���!:�$�r��뿾��Q�h� ��)�Ƣ�g�M[�ll���Sm%��������C�%�铵��xM̰�����~��O�gXV�e��t�y�,%N��-Oa��B��q���E#�tl�@�a�H���δ�D�B���AݑҬ,?�,�������mPj�����||��2��E��AT4�,?yb�p<����ˍ�G{��&{��YC7E^�c�M��^���͢^=�6��ن�[��l�e�]�S܂3�)��'�y6��C2�-�Қ�]$�s����P#˦&
И���������
�֯W{�ԥ~�{ 
/�����O�0�-9�}��O��l�	��"���@���X��^��~���#��1��H�cng�U�骲��딣�k}�RNO��OstV��S��2��f�g�k�.�|������K����l�l��b���dq���R��q >V�jqE������܆F %���6�����&�"�ξîTS��^����<�Xf)��L~����8�e�%�c�,q�i�U?�x�᫨컇�n�w�����hg�Q�(��ֻ��_��jBy��E���]�<�{�$OS�8��ˡ%���K�-��D,����e���Q�'W��=U�$�Y�� �%Ry�F==�"२���|���YH���u���@'�\���g��3�Jhf)���)H�/3���\EGA����;,J�ʭ�Q�"閸A������;���8ӽ"��0o���Ϥ����y�o���c��n���|��ŏD�D�*t� :�I�����(�$H���7�t�l��tK����h>��'_x/L�&L���n��c�2$�ؾL����%���1.��atᷢѱ�(;M�g���򬶋t��fv�+OQ�1e:x2����	-$]b��?,�Pks"*�����x�	j�n���V���;��.65�e'�{���g0�拑R��ƃ�Cite��r�D>�������buƤ:t��~ ADnkzf�s�1_� -hY�C��D��f㜧;��䠆9L^�Qs �ќ����C�(�4$`��k�IX���m��ǽ���ֽ�oz*^S��z��+Db��آQ�������b�Â�[���{o��� ��]O����R=��h��;�eb�t�c*��x�ʆ�¯D��1Ր4��Z�n<�K@�gS���=ڰ��it������,�#ϒ���<NÝR�J��� 5�7�4�e+>bm/10�7�&�h��V�+O�zhTb��׬��H���M
�v��3-�Y��a�S�蟊e�}.$��c#�U懜\�?C*��Rt�n���x����s��2�� ��%��_�����t(h}�	�Bx�E��Щ����_�Y�L֗0���X���'s���F�B��9z��Nǫ���ҌH9Ly^33U�zUTWA8;�5����߾%'�#��9/�A��T�見�̸����[�hO�`t��ܧ1V�_�&���Ht�U�n'�W7�󮑵[��		v/#ɠZݼ|_F��G$8tSH�Q������z �'���R��}U����իz1�^��{�3��E���om�I/���S�^�~�#�2�SS�ZF\��_1�Zt���_�?���������ǀ�=�2��Hr���w��Se!|�+�9㈱�!�y�D���8�@���Ñ ��e*R�V���r��w�sƘ�w��f�'I��M
OB�������%�fv	5�x���Y���j��[�:�pl�qZ�Wq�>�MR-�+c��++���A��p�.�S���f�&�z留M
3^eY��k� ��!�CmہT` a&k�=�}�|m�0�1	� �]��{)um����Mu���S�����)K.��v*�X��n!z�$�+�0������>��5���"�� �L�o��c�)�?l�p\UU֝�y���<N,�y���i�Μ�����V/���hU�լ���)�쵧��r�:�*Ƶ
n3����2'-��I���5^�E`�E�>c���g.T	���B!}���4����t,�Nˌ+R���s�V�Rx<!�0��/`��df���+�Z+��ٝ�[\<��V��^*vwxp�lJRP?��B3N�O1Ovɜ�h��zbyB���V�|�V�b\7* ��*3aT���ޖ���6��T�y�G�=g�"�5�.���s�
��}nA�(�NQY�]�9?F��\ ��E��V�� ���T)C�o��~<����ُ�&u1��Pl_�9Z������T;���M6�Cb�}�<Sf��MQ!���^=�X�;� E�o��n'���F���xq�s1�e���z���N�e���L�FҞ	Nx��CO6�d:�|,�6��A�UJ��_c�i`ʍ�zO_[��]��	G8��=�ɂ�^pe���nS6L����m��H�����U���X0��V����f�.����z�4H�0���5A���(�3q.�{:��׈ُ�n��v���Rp[�9Ǔ$|�<C�JB�~��7b>&��ۢZ�	�2�o�,�!]sK6��㍎��M��ų��F��RR�|:�(+�@=@_~}`a]�Uה���y��s��e<.�(�,�_��#������Rt��=6v���aCҼ*-��l��[r�a$���xre�_b�l�.������E �Q%��N~5���%�Y/Zu%�[\I)	�+�W�����/&�Eۈ_�����]��-��hf�/�k]�6�.M���MN��-�/a�*�J��Jp�� f�f<-����߁��(�~�hP:�t*�0�������07�s:4�` w.�3X%�Jػ���f��/��*G�y�����M�ٻ�&'A~o[�TA��'�$اv�Ӈ�=��3*�s���5$ !H\t�m�c��nnz�كRV��dp�ϞN��W� �K�j��� jJ2�Y1���.��^�()���`���_���DU��w�D����N�pm�l�˛�溿mN�CvJ(ˮp���W4"�m�����Q�i�ң���&!H� �%�Fԭ��������Pɉ,ӞS�V�l�	�}�3��D�1R��Q}ѣ��c&K�A���#@C�������!�t�-,�5�˿�����3�t�b�X�	�@kǾ{�wX=��V9]y�1)y'��V��A���q�S%2M�4��Z4_H,�S�B:�e
��OKlYPǬ3A��e��-����JȎS���ޢG�[���^��5�R?w6S�+E��{�^�*��}[���B+5��3s�Z�V�ӭ �XV��j�52cR�~��`���Pwۈ�����:�Or��R3uʑ��v�,<x%�<���	Z,g��	 �f��B���n|�T�Wj�m׆�i�9B/���#��ѩ~9i}. Q����9�����q�pѳWf��mw2l��c�W(۰��I�6WM�aac��̶k��:��L�����â�"ֶgQwU3�Ր �5��0�N��q�e�5~*o���^F9*!��I����֝$��AT���?8�%Ls��w9r�cF3ۙ�������V�/�"��b4N�;��BSZ�6ۉ�f�N؃"<����]�9�%��Sz�5�(ae���5��s֫*	�O";hi�\t3��̯�*���O����Ny�og@ɳe�Y¬��_�����vn.U��Te��G,Y�w�:�<E���gD.�$:�n�@O��
�[�S�K��W���Oئ�-�ə�?m�����G��\�qZ�
g"��["�{L��^���)�B8�Ɇq�Ԗ�[�Һ.��,�^�%��ŋn�\.��W���vF��?���=d:h���₰��i�D�E�I�]F��?�m�Q����m|���5+�?qҥ�3�A�\ښ�%!xs����C5�i��G.k��/9�b�s��o��u\ԁ�D.Ёw�cz�<!쌓o�O��A	�9�����{x�{M8�7qb88A�y������WD|�Y�}8h��;59E�E�|:	����d�\y��	ɍ��ܯ���M�#N���|���T�'�w����F��n�kb�m��4�Uj�I�R��6�1�<M4�]��~�D�(����jusC~n<�	*jr � ü$O��zVDhf/Sq����a�Ђ�/��Q�%9CR�D����'�@���T��1>;x��Z�<�p��I���H�>.l{�������J�;B֎��$gDr!;��{���NTѯ� ?����1M����$w�J��&�NS���F��U�<-��?km^liWf���{Ǵ�����O���#��c��ܻ?;�J&ox�=�)�]�͸�&�w�?���0�
�:l�>j�Q���U$nv��7�y�gVM䠿�t �R�+����-��^*�k^b�y�����B���f	���)�����ƪc� �?A3�qO,�ƻ/��-��$�
D��f6��d��Qt���	t����;C��K�U���t�k��a"��H
�g���8���^��[&���nnCݿ�����fJ��-�\�~�jś7�f"϶!�W���x��-^�	���I	�!���=����p���T��ɔ�4��,�D�_z�|_0b��u��H��D�d7�p.o��v�j���C��6C��U'�=�w끝N�⡵��������y�SΪwd߲��(�+,b���7:�P��ȉ��A�Ud�n������&<�7e��1 -�/��m����-��;��dX1lk����8dHJ�@��j�������j�,�b�>\U�=ya�� 5�E�}����~�NǠs�-�o`1���X�mH��e�g �;:��ʲ�o��^�Xk�����-?�RE=�X�OQ��>A�O���E�������y�/	*��j��[��g�@�<����$���%"^�����]:0aq˰���-�*����{��F$�,�ZZ�)���`3b�O��T�PG�AK���	�O������L�X��r�	i��Ǽ X�xI�7�˞��an�,���W��=_tyݱC|ti��/V��������%��Qu@���w<���v�4��Z��,V�c�9��?� ��_d�bfC}s����2�w��� )N�^�Uƅʊ�w����f�0ทב��* p��9��d)��:��}��Iڣq�{��k{��M+54��;n�/�$y?��8|�|��l)�M�=]̷.��g+�󵠾�##h��e��#۾Og��(<�8j/��s�ܭ���T˸J�cs�����R��Xp���::'��Ua�/�K�Tx�v��\��<�c'�r�~�o���~��]���]�(��wŠ�h��y����}@YO�/]�?jI먨�qGf��|��u����;b部~L���	o>raB�
���}"�=)�=�Y�k��;Z�x/���4]3P'�c8ݣ���^C�0�O���U���A\^���ԫgd!=Z�+��Z��KB�~��.��)��brxY@�� ����\��S�ct�0�ԉ-G�r2U�dl�z	�0J�u9�����D�)W0E5˶�lB��� �ۗ�6�};`���N�H>E.���6����-ΐ��I�]�2�F�m�_.��>	n���	�͗�S���'�^��Ir��\~ �H2�A�.LE-��`��T��S����i3SX>��D��kЎ������S�K�T���AO����a$�%lZ�&C��}�:ɼT��0��=AJ>�\'�דkƏ�Z�D<:��o/C\�����l��%{��<KvW��.2�7�6z[�in�O�&A�=��.&�� C<ň̈�����u\��)L��v�Y��v�6�BLYr�Z�H��O��n�hE:>�A��?�9��)����1�G]��(�l����yv_(��}+W�,��:|��a�׍�!���Ueŉ*o�@ÐT��WY5�`��_�8=�׏a�o�F�zZ�nwa|h_}�6���À<{D,a���U�ag���0�ˮ�!�g���~�snd����ҼR9vVqD�b���Y���}e`N�@���L,�o/�h�)����P�No�B�,^C5߮z���(�)l��G��e&�'#���~	�T�,��Ķ��&�'�s�N�k��`ů�I����B1c�_�t��m��4������3$�k���*�<>���la#I��H#��fk��� �{� L}Q!�C���Q�͸6��.���V���J��1N����-9��Y.��ny����J��;����
F�&����mȨG'�f�	<�XR���0֞�3� ��E�X��Wv=*�J+Y�#���"�`%�y�/���0�D'�g7�&�;4�s�Ҏ�۸�/��Y����>sȝ+�n�d������k�|9��ϱ�#`ø��_R���T��v�rz�?�S̰uJ���h �I�����6��{��>�%Igǆi��6��\���5w�w��P�9ґ�)�w!����v�����%�ܖ�乲^[��9�-�Q~�)��]�_��Q�+q���5r��C��YT��H���lKh!}-�Nu���������N����U��u�͙�p|�(�]@�}u�����N��pCs���L���Jr����1�-�oo�źDa��j̿���W�����5�|�Χ�\�Ӕ��mt���L�~lw+�SP �+�3~��eͺ/�0�,WV����H.�7ϣ�r#S�%��b�KC:���_���Pr�S�W�2ZW�Z^B8�Z��kʶӗi$
���b��k�����r�����O���7�V�<{r}�4��^�uLtغ��t����gf?�L���z��I����*V�k���ߠ]&w�����?^�U��xQ{��������(�6�XXn�J���}.�I~U��V�6�i]�u�Y#��z����E��Rx}2�/~�jΑT�\!��|'����u�m�;����"��F["�O�\kr�֚��؇�?�$a&m�������$����X����~����P�/����-.�g;�d�?(*D���bsHki˛5��+/��������4�.Ql��`�8��~�9���w0�Mj��W��Ր&D��rw<�������":"f��}Z�!n�i:?�\T\8jY����eM:R2�����5'�P��Y_A�l��A^7y�y�\�u:޾t66%�+v���3���C|�>�wUo�ml��a����>W��������T�V��Ý[
��b�I�Í���a*�lL���D�}i�.~��T�Q����ľ�u`
0�5Ї�?���WxgXo�ǊY�����L�󹫯u>Á$[6�?��F��yGH�F-�>�5�7��Bg���mM�ק҈
�c�۽k���X#GHYR�"xW��:Dݨ�7��)6���]EtU�g�هwE
�����ѐ����r��R�NT���g��m�-9�]��T���{
����h�+�w�2g6f�,�Ӫ�oh\��I�u�Ԭ�>�u�-{�z�|N;�"����Z ��w���3�ĸ�>�&"l��'
�o{4�,~$��OnT�o{Y��ېHa&�-���?o��VtVк��&���H�3�x�-���(	=A��8Dتk}���q)/Â^�
��1�o��,���e�J��+>�d4�\��� �QWN8���W����&�Hg$��n�a�盢UcA�u�&�`7/�V�B�L"0?Q���N�ڸV(#h�&�i&��u�˕��+>_RE����B|����r#��ݎ٢����������%�#O5��S�.�OV��[�P(ms̀��A��:���|����t��[�'$�2+c��� �i�j\>��χߖ։
�V´�T9�w�%���Iݮ/j��L`_x]�AJ��h����9h�A���z���F��X_v_6����6����<�BE[:�RD�&��R���D"�]�z�s�TJ#|'-��xq��޻5ʔ�e����+�|i7�w�#<^0J;W��Mm���R^��j���[!���\6G�mH��[ڶ�������o�e
��x�_/�6x����U)5{<�}E�h�EI�X�/�`xh�6�$�����k��b�4��s���K����q&���-s���3�����Y����ldg���"�H��m����QErx�������*�������ʯQ���k1�m06�������Q��n𗱈��n2e[�?S?�T��^Z��%.����x	|	'���+'>�f_��H�/���7[$�'�zK�4!�����&���<��|��T��d�K���^i�� }qO�����5����f���ȇE����Z��ͧ�vv�A}�������8W�&J�r�?c�f^�AMX[��lO �K@��B�QΔYkQ�2<)~[���m�+
B%�j�2�L������7Q����~��fOK�Î�����7$��2H%X-:��������gP�;�{�2��C�
u��~v�hMG�#X/A�\��3�@�j�	-�x�+;�m��M������qT&�ie��1�!��VA6�V-����0���n�zA���|��-�2�)��Nҹ����K:��葖�N��{��W�����%�CDTx�{5vE_2�bs�d���^�S��Ψ��v$n�6c�J��
f艮���>���)�k[��4�ʘ�pd��$:Jw3��$p$�R�w/P{��F�ﻷV�����c��o]�JD����9낢�+��
V���×ژ�2�'Զ^ƍ�����	l
	U�Kw�Ft���#�Vsn�Nq�}}���~���m2��\S�E^��do�� z�Hv�b��?�p��M��$��K%\+]c8&M4�z��4O�G�'R���(��t��s#���H_*���mY����|<���F~����;Q�#�WlwZ�a�L�v�0ߨgiU9`[�c��m����i,�k�4'��!2Or	�_�mT�,��1�.�Sk�*�%�P-C�2���!���&�6��Q�b��5�֙�aw醂 �n&�K�[�6����x��+o��*�9ޭ{]6��;4����W6�h�1X0SvC'��@�^q��bI<c�N��5�cZ|9@L�+�0�
&�X	� �Ȫ)�-,y֛�5��p[)��Ï��c���$�G�l��~'�OC�x�>�����M2<o���E'�6��Y5
^f�x@�����	�;§�0v���7�֬�bpgQ�	�a&qpY�f��A�9�+'��f�����s�˳�Q�������'�Ft�~�-�k�|����Q][��"���Ū�2P��74E����^\��Kx�5�����3��yJ��D9P]6��n���2���|����M"�om�m'*�1�@/�_^7ܷ�@[������F��!QEU�E5�Fk���hn��n�������El�0l�Nj�IU��-ʯ�)Xb(͓R����Ѯ۫�B��A�;��� ��:�����P��o��36^��:O"2*Į�1l��&�ŏh��N��-�����~hj�V����H��J��vޞSP�L{��|d���e3�4C�P�BU]�n��Y����4j���>�m���#:���/��7<�µ���+�+�(�[8';�w�f"�]I����(vE�2��2���9�jF錜[l���/��!c�
{�9o�<�e�
_zy���u(��9���j<
��z����q+]Ƅy��4�ݏG�O�M����0j���fSڸ��\����ȣEtp�囦�}y�Ɗ��Nb\� 'rg���͸ɿ �����!�F��7����1�j�@��Y3�q�eV��.���>��@����L)�>#AK4ٞb�1��CF^d$�z+��劫j!͢wV�V[�9Ѹ��T}��������".�Z�C~rn:RD���"�pb\���D-
^�����v��t��a%z�t��=����Qi�=��Q$M��El�G_{�h����%} �m3j���m>h �I����S��v��+)9�5�j!�i���>F�������0����k8�	�BL�Ab�l>�.�u��3�g=vg��\��й��hc���/��z����K���s�W����`ը�Q�"S�0Wi��u���M����L��k>Q��BqȻB�W�	�au@����"7rϛ�nh�%Eͽ�+�6oX���]�ŋ�:�g��m2��t���c.��\�����|�ʗ#5qs��i}T������zG|���+��_Ƥ���n�~����?����t���7��C�k�ok>X�3r�V��ʹ�]~�X�P��Lv�ܜN��4ag'�%���G���2�n�}*=
�^~��w�J@C�r�n*Y��U�<�ج6�ۉf����^^�8T���XM��JB*<�$K�=�k�R3B�;�*�eJ�G�\�A'y]x8+l��r*bҹ��D���NH���Dm���q��%p�(���� ��?R��� �Ax:,#����d�M�	iڊ�|���a[пp�_7
����mwT(�ӗxwb��h�8(�<J��rn;|S�{���p�0��ac�G�����Q�(�7�M�W�w�m�yVo��8a�~���y��)<����HbgFr�	 ��z6�Cr)1-�R�sb;;^����]��me���Q7����RȀ?�)8=*��D�
!�����ξ�P�n�ѯ�Ĕ�rsy�����~��V,����')�y�GtTt?�V:�`���uu�:>Qͽ@��]Iw⯣[�1Xc�|�Q���6�����2E-'��|��ɵ�$6���l���R����f�"4��}w�I��Y��z"�j{�U���O��Ϋ�}�1��m�ɞ�El(7�{�w�i&"�Z���:Fa�5�V����\�i j�R�ρ1�剀�l�lw��$�U�^7��g$Kž�����jŦ���&��Op����;��� t�����U[�?:�W�x�we���=AI���DMK�7�򘱦9�Ff�-�/u�	�!�:�����W w�C�Y�k�d�%:=7��^w!�aɃ;�w�ȍ���;Vו�3��n��W�<L�mW�j��Q�]�j�%)
�E�m�j�<n�ƽ�Sz�;u)���sv���+��͒v ��D����x�N�ug���d�Y��ry�p�WrĦ��L�@��9��l꽁�r�3�y2�.�c�k�#0t�4��D��c4��Mt�5���Y�?�yi�:�h�d���?�b�Z�"]�/"W|��z���s~���#����������c�Ƭ��b�Q�0��,��u ��M��ΪFEX;x��X�i�?l�h�_�ލ��8͆0 �S��y��/�H�f��l�
���?�ƏMN����	u��~��QǙ5[�s���)2%��s-z=/9)����L.��]"Y�v���<�g��a��5���|��PEx��1�%�eL�^~�R��/�W�0�K��zM�r}opVۀ�
��̪��Hi��:w�8?�`eB�Oi8r|���j�ݭ�ĺ�����J^FB�i��E�l+�͜1�<�>-�9�u���ڳ�:6*�+P�_��nS����N�^��&��M�Ps[���������$�p]�&o��xL���P32�>�>�8�S%b?��KG����7��Lj/�5�-L2��M�ʋ��vgft�MJ�?o���ʈ}{r���	iP����2U�T�� o�(��3���u97V�z����\�m�| ��t�.D�h��G��t6���ՠ_ccaY8N��`�o@���� �WR����xx�)1��Nݍv���=*���a�-_��C��
�i���M�]�N*�?1�))��i�[N�'l�#�T�$��V�,I��l$�4��^CAp�^t���׎��K�n�΋K���6�D�c���F'�9֗�b��m�&�;��(��n��Ю=�R��m�VR���A��*9b���#{�P#J����>"#�q�<��s����=�U�CW�)��g/���!y�	"�9�8r�-t`���Eܐx��cWL5�7�7S���ȴP��M��/���JY���:���w;�5͊c�?N�V8��@�3)��чO�fU���N�k�U��{l��q����
��&��FA��1��(�Ts�C����{5��(p!��j��FЂ�͠܈7~^wXN�RB��֗�t��w	�Nێ
���K��d�E��M��H��� �E�Q$��n�U��*`��7(�����>吏�z��^��!����x6F�xY � B~��t�e���,��� �$vmBn5n��*�Ŧ�O�tX�v����@����x��T�׍7���`Y��z���_c{|q���A�����˕�gW�&�>���T�8�r4� �����a�${�� ��먴��aP�:�fH�~5�È��'�Dx6�������˫�H�V�� *A�/��<�];#��r*�7�m�"xmT�l�mI�d+���_n������2p�64f�UH[魸Rhl�	9�m6~�
)Ù��hA�;��k�=�����������p�3��p����<^\/��#�
f�c�.�A�i�0�,]I
𞰈N�m�^��YDvh�E%�BS^��p�+�7ӹxJ�n==�q�F�VS�Y�w�2���f�c*-��QɆ��{����3@��8�p���	oƗ�@��$��Ξ�9�_�:����� ���n8T�t�bT��qz㆕��/��-�:7:��'"Aɿ�F�+1\4�|#�e-�	1�K��c?��\^��@і���X�ó�EeZqҾ��^p���:�[�"$�e��h�O���ȝ��Y�)~ L�D"n�B������?�H�1�*K�Ǿ)�ob�,����Q,ɞc�Y�Q�CV�!�FԲLN� P������	\�5;@����s(�/����5�%Cо7�C���TO�ۀ&��o���Ű�(�&c.����8�$��)��7o�����<%Y����5��L���?�Q�J��= }�>b/�S5�{F�Y��\�ؕ�u�� �pB1o��+]�k):���6��^���C�{"!3{�5�h��#�KPԟ���U�Igǂ�*Fr7^nR6-��=*�w�٣'R�Ok1�;��6��G=/1Cx`�xE�j�������壯����oȷ����
Y_z�xa�ri�!��7wט���Hח��ۛ��b�Bt����d����:��[�8��>�U!�^�ׅ4�Z�G����ۀ	�t�:�C������Xzj�I�Kq.Zt��ތ~ev,���rE�� ɨ0��Y�u%�����8�b�����{�t%�;��Y�������&���B&��$u%�9$�vI�M����[fě��P��z�˾/�\I�{�݊��k���	ů�n�����;�b��(,m�x+`%q�Y�~_��`��0�����`t��Z���A��y��O���f!�|d�.��U?�D���'�����l��9����V4)��>�2�F�mM~s��y6'0N���^�mPG�;2P$������Մ�����8lW��K�u�����%�4�kM>�X��x(���&B���S��%��TB��%$&K"�.�]Ǿ3��=eI�>F�(���{���������|��8��s��u]�u��-����\�jP�Y�˒!�`�!��rM��)�5h�p�(r��h#b�����pY�Bԩ��7 �fgvx�Q��s�Sbi�?P�R�vu���!BM�*˼�M�a�5�m�}���-ZS�
�Z��#����(R��z������=Iú�Ie{Rۼ��KQM�$wp�.��p_�a�K��=[GZ�a�e�!(u��z����	0h�w9wٽ���Z�H����ڤm}�C�n)�]˺����:���;���ф���O�J&O:��Q��*8A�´�[_&F>Y�s,bg`���9�~��vi�s�ίI��x����0���`��)Q\�Ԕ�:���{��F&$�j+ ��ځ�,roSտhG�_b>��G>G��IRH�i��KM�2�U���� ��X�8iQ��O���������)*wY��B��I�	����X�]TP������bl{#�|-�d����!uqz�Mj&	��AjbH�Y�FӒ&�U-in����KfQ϶�/\�Y��W�E>��
�y�#,�"+-�� �Mv�q�ޅ�vYa�>Ch3�$�� �Mp���h>9]��t]�8���,�D蝐R��-]%�A~2�������&���
G皐�儃��)���Ȭ�Iq�@L��E� 먓)м��K�QE��C�K��e���a�M��׭JNZ�/�;��MI�~����۳PpB����E�m5D������6U�b���|sHp��\)�c�'C�}�cOhP�H3��Q�ѫd�*y`PW%����h<z�n��p������ȑkgy����d@����-�>�ہ�`�Y��ω�^�vsq�	��ᓐ�
�_n4+����q���e�eu(F�z`�(��P�#Ċ!��S^�2�=/Ȩ j䁹�5�	�r��ǎpƥ��ۚJ�cH׃���J����� �7vq5����I�i��Eħ���o�ȼ��r2���ctĨ�@Y�����y��Yzp�yc2�w�gI�6�<A��� ��{������#������I�E�@�s���_7�nu)�	z��"���7���&w�Ñ��%�'���}k��J����~D�'(3��l�L�5u����W��Q���%���0��#��0x�o8�e�f�݁�#�ڴ)�:V�ҝ�_�?�+��%q�d�T��v5 x�ʰ���ꈮH F�ɶ���k�ί�����#,���7z
k�ȱ��^�ۙ��I6[
�*Y(�T���7Y�K�e�B!�N��`E������~dXs���{��ЊW���E�7o���հ��Kv�A�r�l�1�:?�L�t$�3M����G���QQ�W���\6\�ï5�|�B�]+	�����S�6���_o�,�D�1�2���-t���_AQ���(���} ?O�0Ъ��njN��;�keB٠<'�Kq��Ƶ��b��|
Ւ)\��(����#�K�;h�+�#
.]L&U���[�CBt��$����;�
!A/�w�V��T�eȠt��BnȤ��*��/lJ�D�ѹz�0戈&�c{8p%2��c�#�R�-�k6%�n�Ǧ'�\e�CY D�H��9<r*E�R�i;�>�����{@\�z�4�#���t�[F�b�A�O��s48p.�qً�bH	b
F����Oe��Yk85��v�a��f�]0q�Y=�M��-��A@7�����W� u]�9���
�Ļ@=�z'�`���9�Ȁ�oƍJ]jy�S���n[�ej�[T���>�-E%��C�(�-��)�U�F�4���x�:����V_��֎�ǣ<��W~v?���i�nȣ��2��*(��o�`��&ȗK�"�Um��Q�%�Ju���5$�e�j<-*�;㴉8�+������L,H�@�<
���$�Ў����^�}aX�(�Aש���㵁��Y����ͼ�/�9��!�\=�B*��5H"u|�z��o$g~N�T�S�?��F=	���
 �~c�P��*��vȾ@���PJp)jX�V��K��x.j���$\nXiR�W�҇���tן��3�D�9
�:6�2[���@�^���h�^�@�K�a�[�p�6�O���;	o@��� �w	�����$��V�4��r�}]�yg@.z�M�e&��w"Ѱ!�����A0� 07 �=��{z��� s�u�*�����Gع.g�|U[N�q5���B����:�K���]q*�9��u�}�'"z���\L��v@E1�o�	u�ܘ�����;<�},��Sb��@���r���%\0����w��ZZ����Y�(�Z�vw*���(�dSz��9�x�RAٸE`H�1�x�ݪ+K�Zؼ�,OaN��L��-`!��FOL��l�џ-�';)v}\�I_�=ҏq�j�f�x�P����DdU�t9"Ɔ ��N�xS�����2���?]�t�$��%��|��U�+W����4�#"6��L���,���>X�����0�k���Y��z	Uh�+&�2����f.jrF{�Xo��"��x��ۜ�7T�� ٩<�lRAzu0I���9��zP�VNȵ��P�t�:ӵs���ig�1������{_K��)��$���0�d�l�����n�9��*�/�q�E[A
;�Kk:�۬ѸДc���ӑ��P�ka�V�]ӯ7*�Wb�RO��󺎤`>+�}�-/�C�ɕ����#� YDeR��润�C��5ȏ|ҙ�n�=(g����,|�%L�����!�۬I(LJ�E9�k�X;���K9����I� @G����x�E���p��!@�ˣe]8�\xx��~/nxR�i7!>yTb0�v��$�;�v�>�\N���x�}���q@�R�nG��`U�Έj���߷�_��{��JP�PP���f(�ꯔ3����qw��x������޵��:jH`N�=I��΄&�-`C�"q�t�8���W�Y�{U�M,{l�H�[-�b�_Z�f��]���b/�'X��d|w����7�B��G�6J�s��ݩuy,��&�,��q�'Z�9���R��!��W�t�M~tKŝ�o�*A�����<<ZHF�PM�*|�yb��}��r��%H�\�	!�"K�C���r�v�əh�L�"_��G�޾Qq7��`��}�S�����^���䎟`��V�X=�3 ��(k!z5�O��k�I���:W�U��4���v�a���w�(�,��Ke�,���7�R��,�;�fu����~s�/�q2S*W�� �b��/��]) �(Q�#���KԪ��R�[&�U�lEC���.�]�������!ً�w�a<1��:����Si��/J4]X��U���������c���鏝 �;0�����<k�lL����_�q��H�۸�����dc����|��_�W��_��{��'�T�:���!W�XfA,�@�#�q+�e��aܤ?)B��/F�[i�!����0���)�p���re���ڿ�0�Hbm����ձ���Q��s,td��Z?���e���¶�:MD���g���!�ض�:��<
�Tb�E�j�'Kj�е�i+z� )��Y��bu2a� к?H�Zǫ���{JQ%+�� r`�B7v�%mo�_9�|qG����Ư��U�#�
�ؔ���(ר�Ð7ֈC`������_��^�T�E�bD�v��:܅�J�G�3�PE�N�cq1�m�D ��q�E��C�+~Nڏy�2��t8�eEi`K�z3�͎�d@��&Ϥ��D�;	��2���͕�U�R�����e3h�w=>r�e��Фԏ�pe쵋��]-F/h�^k.A�r�I������X&�>&K��ċ�I��.G;y��z�H�M�������>�e'��@�WF���ǲr�ݨ3��r�^��v��RŇ���%�S�Z.Z���m�9@!�r��4�'R����o��W�v�6�;�t1�����a�6�0�v����~@�����.g����3�r�v��@E*[ƃ�ߔ,!��w�xٶe��c�kl�k �%x�5��>�_�ŭ�tc�>M>�� ���*��6! �<���}@I}U+T �V�v4��>	����H�?	+vڐ���I>���������^X�!�&(^��ސjn�-��"� ��0ӽ �r?��]��
�@�mq�gۨ׺e�P�/B"Q]!�{��g��2��h��3T�bz+��s͌&���u��Q������5��Pt�g���=�\�{jn�b��a�y��w~0)��a���vá>���NM'���Zs�9(N��b��|�m�D7����D
v۵�Rz���p�����41i~6o�܋i�J�7�c�7�u���SFU�V/�λ#�Y��r&�O�mq>�%��� ����ˮ���>��w���6�n�=C��"T������K#�&G��`�O��ll{1����Mb�@}i$�7�ˌ�;�ϳ^EI=;��b���VG�}�[Shp5g@�ʆ�Z�J7:DSB�,�6]�޲w��~�Dw���>�ˡ�d[Jk�(�(#�(�Y�-����}�Ǩ���򠭁9�Ӄ4D����_���~|�L!����׍ K��5=/�E�_�ܺ����I����G�D�s�b:V>�q��l�5Y��v��%Ҿ���x����Պ̕+W-E�A�6/L�I��Of5OI:w1Yߓ�ãI��i|�M�{��Kw:���Z�Sc闰�=���!�%�wT�;u�k�p�H����|H�uIG��~�
G�.VQ�;���<X�FG*�/�]53�`Uέ�Y�Qv5��d��:�?2d�ϋC6�֜�j}��wj</D�~t�!��܁���@A�f#���t}�'˥�&�-�S!�mo���е�q:|�Ĝ!B�.��2$1i���_�����1��稒��sl�Mf|� ���.������h^j�4��4�	^�0���4f�a5 �I���ؽ�F����4���S����NW�h�K}�������(L�m��g��	��Wi��0��'$�~���6D��󸢤'܅��J���������w	�1x��C�^= <9`ɵ���4ɠ4�%��/!��jA���!œaz1!�;!]�M`��&�O��T�_1��"�������F��~@a��}�g���óv�bg��ݺ"�m��� ʠ�#I������I�-9&�Op8_��n��p({��l[�����u��s#|dq:%׳j_�����$
U�������L��Ў͔�0�[X��^��O��؅c��z��q��6����#8!��D�+ �;6�O�e�7���{�~�,O�W���f�h�X)�`p��b�qڔ��FY��Y�,���z7��������T�~؊Չu�7����'ҙ�Y�%I�؈	v&��*�MS�PwXgq_��Cg�`��	�u#Sh��W�y� X)�Jd��b�ҡueW[r'�?k�%d�s�e��*��X� ��6����א��[��:A9jR`���s
�$�ɕ���aNMk1y_*3�������9�z*�]5�u���0�jV��3��^�9&��b�*�Ӥ )֟��K��2�'F�6�@�����s5 �Ӏ8Ю��%Z#��
d���<=U�����x�[��V����w���q������g�Oe���]�r(DW�7\l r�!�0y�&��㚝q*�k��o���O�K�.H��=?%��_Β�׍Le�`�r��&�r����/��wP�3���9|�L��Qv�pI]�v+0����7���`�օ��?wΠ"���Kw;*��L �9+ѣBK�:��Lf�=f�]�#�A*�A��f��	B���>ѠB�׹>]z=���o�S*�މ��BB�g���~X�?�	w�����0`��&�	��@IH���G�^�T�0�����k��Z}4!*�J�C2*yt[a���h6&�} t��#�#�ɰ��s��H����?����P�WŔ����a��ضN����XFS�� �����Wk��\�oz�KX ��sMdS��I�����P��t+�c��ʌ-�Zҵ��牤޿�q�|H��%!�HpM���q�"v��{�΀:.S��/��5�K��ڢ�J��(���Dgb�� ��:��ju'�4�(��Nog I8� /���~9v���gj�mo>���@2�4o�C?SjI1B���Wwu)�A�(N�D�Y�ܭ�r͈�m��hZ<w9푡ޓsE8`S�o�.j><��J�4CtX������G�e�G�\��t�[:�34p
�	�vs����sk�K%?&��/u��-�Jf���F��V�k1A��4[C:KT�]�un�wT��t�#��I�PWp������� qxk]��Sj�;�\Y�����&����LDB���4�H���\�Çr�l��@�;�% �g|i�ۚ~�K��l�
�e��~]zij`{��+oLK�;$�{�9�1.\��f������g�����3�+y�����xh"č����Ɋw$������O�=x�����-;Wkr�VT�Y�$<��S�JQ��)�l�z ҩS��S�G�9��l����OB��Q���߶Ȇ���~}0ݠ.�9*���9$�%�w�ye�s��Kxc,�L���0!���X'qL����r�~��L�@�������Y�Ko�x
��%?=�	4��}G"��nv:��މ�H����K0F���0G\b��lex"�H�.�-�@�\!t9NN���Q��Z�'�M�ӛ���L+� ]~���!j�}J��w���2�r�D�Ų�t	�SېK�raRꝐ@����إ¾+��h~7T�O� BMq�'��Z��/����$|r?)��j�_#[�!e�X�}��![�
���hY�e��� ��`�L�t���I��Ւ$P�oG^ay�~�s�$����L:�V��x�����tV��k�"3�� ["?���r��_�*��G���N23�)�Ӗ�&�����`���q{L�.�+պɉ����A���?%��6 ��*[�y����PX��3?W?�������4�<��"��{	G�dS,���6��x�B���	��U+QH��Z��0¸���P����evԨ!PQ���sq'�0����%����Ƕy̑_�˩��l�V̺K7h!�Y����u���qC�a�[�b�x}A��ȱ^&�`c�̞l��۳�PG3�g^o1���hcZ�5D�b�z�jC�Rox����R��.�\��i����s ��U*P�6*�:�~Ҟ?��Hu��,I_�q�2�ҰW=�h2�Su�����[N��V��������-�vqm��v-2E�d�����Y����M�0S�S�:�E
��戥%u�<��J_$�prn�l�^���E�=F@kg����Uy��<�N����G�7 ����B��;Q�s4 �PsuMǹ�Q^;?�ˈ�h�#�D�O2G��}OQ���&�z�x���{�t7k?����w�nU|��7?�P�.��)+[��@JC�6Ҥ^,^d1��V���E�K��:�� ����>Zf���D���=ȩ��M�0�~�s(�{�;l�֤����>�X�5�G�v��w��-�t�*B5����d�F�e�A�b�?�̹�1R0��"E�w��b�&��,�����R~*<�A���ܪN�y�:� $f����ͳ��65�Hg��}է�K�r$�E�;5@L��P�IV�;�� 2C%�D�튚O|�0b��IÇb q�X���<$�<��¤��.�`p1��j�/���\�w���L?����
�r�#��<��i���ܗB���5ep�V�"$Pℝ�]|E���c�.��MЦi�ɸ^�Z�b2����4���N����19�뺧�V�����^�4G�ju�B�h�!��Q�R�9My��=�h��6kv�x"������-K�r�G�]ޫұ�\�����
d�R��� w+@�N���#rdٮ=�����K�?u����,�&_�2у{ׇ��&{ԉ�_�{u�݃X�fq�4���<Q����(��Û�!=f��xmK�3^T�z���nJ�6x��%,�H���hQ����w ��&ů|m�����W�޶QA�3%�Ɩ����LPCR{�s���yX8�5�D�W����/M�]�z>}�@p`���r��ǛZ�Os�X������P�� ]e����v���u��B����[���GhO��x&�mA�h���
?��ΐ@������[��(��FGJ�Pҍy"%ƕ;��1La7��6e�~��J���`���2'�WCF<��F�?.gҤ�dqa���֧�N�mZ��t6nW�{Q����!�վ�5���>�Ӈ�'%��9���𯬋��F� ߞ�:���rz^2��F�,����_���!ڿ��a�h�Z����z9+棺�oC�}��^v���;m�O�D���ݟ��Ke[S�it2A�	��x�0G��q]�	�|sA���4Ad5��u���8��k�<�]��i-�9x��]� ܺb��(�(L�و�T�9r���:�Y�q�'
3;��-���]PIƺ��%տ�2kw���ٔ��8y`��]b�8�=�.h��_G�${��ƢoG�__��S���L��+
-�0?3.��zq���\�(�=.P&^wa][�����׼q��r ;2�Gذhd�!����@]P���go׍f�Op����[�fHC-"��8��SQ���Q�.�Զ�@rA9c�4c2����$�`��u����ز��A���}�gI.+][0�t']�P��$-������2����B���m:FB+��/@rIF'�Af��ܫ�ӻ��h]��+�#�l$i���;�x�oN�# �pN��*z�IQw���v[\�I�d0�-E�ή�N��UmL��t�6�C\;^�?��T���8�����_P�9�5@��^�lf�L��!��
�Ec���(�pd�s��ަ��� G^Ua�,�'Ό֪�?z���^�L��.�"��waT~� ׋�hS��ge@B|�؉�]�z�nE��d׏̝5�����a�H"j�.���=�sͧ$) T��Z;>�=�A�������oZ��TD�q�mJ�m[�����]����_�"x��{����� �f*�qٻ�R;A����G�ƉT����x���F2%��߼w�|�M���w���:��?"���׻���fXܰ_M���u�~�+1j1��"l.h��_�0�-���s�Y�`\db86�X�J�d\�ZZ���c��4)�X������)��;��a�o�)xD9Sz�@�
��n,�de�H�ֿ�ڽ{U��աe�C�o6e�l�+S����w�/v��ǐ4�;)z�o��V.���ܙ[�J/E�m<tr�\mb�Oy���y5h!(m������x��jH�3�޼L_�.h`�v(\��jG�U�Tw��18�����Y�DOq�����8ϡe-h����]�Gc2WJ��˟49��]�˒�������@���L��CSj�yJ�ltӧ%dJB|o}���֖���qǪw�?Hb��yM���-�p8d�b@V�
��� ���L�z6�_lPup����V����5��V���(L�]kP�4�p�LZƇ���\�=,��)�3�MB[�Xn���:�_cT�C��@X{�#+}��O0���9�wx]����a���A?�G�­��b���!f�߸����v�9�#����"N�]}����N���̝x��h�AM��O<��z��O"�Y����]#O�M�0߳_�7��a4�S��5��k����t�_'S�������B<@�?YɎ��
Zҫi�ز�AE!�_ѻ��mVᥗ�՗FnD:��:��=n��/1��. `�P�ZǓI\��"���<�H�oȕ��ҭ|6�!�̏vl�Zǐ��R�'[=�a����:�9 ��3��8��ӯ�?	/�z�~ ��F��W��������[�Az�i���s��J�|C]�Zgj}O@ao��ݬs�#<=��4�)u����˃E�iiBiZb�f��|���6${���Lf�X���&�!�TݕY��N�\5�z:('&_RC��]l��9��q䫤��z���1�P�]��Z ���	�.%���dOQ�;�?j���M�^l󏕎�̊x���2v2lp� y�YXS|��}��g~���)E��O��ǿJQ��V2錄f���h��>�l�����b�u�ëF��������l�ߴ���f*�a�}�V>z�.�G�Қ~?^g@`�qI;��~1�7�_�?��%��][���	��v W�FH鉽,���e�}Ϗ�kF��3��_���ib�NM�y�9U����0����:�CrQ�*��I�$�8�� +w/*���5I�b|�J�l8=��2�3��'}�5�rY��m4���E/�)�z����o<�=�w"_�e����$����5���QY�`��eyOש��]e1�1���%��t�zq3��聂��PݯK�sv�K�&�.K���Ų���w�$�U�N�zg��Y#w��Сe�̟9��,
��n�葷h�$��?Dˬ�{G��������g��T�.���T���-@k���z
B���q�;PK'��@�4~EoZp�E�I��w�Ti����3�p�����T8+\�y����h
2?��F�slYKY��K?H��ɣ��w.�Vi���S���*ޞc?eG�[�H���-=�5S�v��/ӛ��[La���ɏ7��Ǐ�5k�D|AZ�x�%.0�L���t�}xjo:�`Slm�k'g���\��|��^�V�y_J���8$i�j	
��5�ںAF��m��� �s��{k+�Jֽt�l[��ۅ��~��u@w��띯$��d�UO	1�у^DIo���E4
$%^ϕ�������j5/d��!��M���F��ФMq8�pH~|纪�7��k���rh�W4�� IL��7*4s����];��Y�X�O�F$.�EX2�j�<��H�V��+Dc/��=�"�z� O?,~\,<S�����mݠ�V��a��
X��ȿUW���	f�5;ٳ�� �d�:��ë���"��t�˜�^����aB܅�TăE��+Ԑ5"����*Ҷ�*�!Y���?"�&K���C�Pk�
4��f˽%r�.pD�0��H���̕�}C5��l�|��������� k�h-�;�}ۧ�V��'�H;m)A�BJ��$q���>95��)��k�U-`��Ei�������+8Xǻ���?�rv!_�%)���``�|�Ǖ�Z���lR�޸y_ �o���������<c��dXs�q���C���m����Nj=&t�����YeĕZv,�hͤ�`7�9o�
@�>z����O���޸��!H>��\Q�e�$��<�@,���dL�灳4ܖJ.�r+���#�-���CqZnB\k~�vxto�ALY�s���i�j����}�5�r���j�U�:�~�IW�6��� ���Q�lx��J[췢.A��vc_�I�Q�&�K'�Gao�����"D� �!��5�CZ?`&�e���Ґ�6s�V[�=2��5������l����~�����)��h-�t��Tt���,�L6�t��+/R�0Lf��u>m�{�Z�?�t���vz����fT��̆�2'��"��kJ��9�K{�
�m��3�]~<R&��K���(���Ź6uY]���2����x0��ű�i��Ki��Te<.k��K��M�e@�^c�7��fr���?��#�}�$yK���Oy���|/�#΀!�Vb���*۲�8K�i3���T_b��@�����9G�I�)Jq��֑0�1��z�aK�>���nk�8��ZBKbm�>8
� �w����1������yh(��m��H��K�W���� ���~?�y���˳F ��%Lq:th�[&W��)wt!����r��:�!�H�%��{<}mg��ӓk��6\��z4�j���ł��Yt��0U�t���O�7�hfu7��8ho�a����a�Z���]��V�M�s�o�qt�A\��5������[p_�*/���}ߔ��͎�UD�8��)�\q�zm������Tu��oU>RJ�Q�P=9s��3m@�?�вp�uV�����6�m6����q�qW��i+b�^.�q�cܻ�Q/<t�}������t��h��î+W��~JX�d���ӃG��Z���|%��e�!4j^<=~'��\�����NF�$w�=Z�2�RN��֤������2�/��W�`n>����$����z�K�
]m�aƿ#�Ju�1]CA��R�}2���a����Aȍ�������&n�.���^�.���zK�?����d��7� m6��ILG�L�}P����/L��h��,QI;
`�ω����6�'����4��h���=k���;Bݗ�R���uee\�x:W.�G�� m�o�\0�8*����M�HWS�h[�%)\Acy0kEM�5G+��WU�/�#~�S�+y=}��f4�1:��2�����>���b��8��l;:���fsX�,�_�Z�>,�(��	��a� .��%�OoMp_�:���k��t�\ ��Ơ��vf�w���B�QɒoĆ<"�!�c"Q�� @�=��x��W�p׷bɒi�S$[M�8	^���G�ۉ[�4�{	��߷�m��fSVI�Ã�������hL9H�
�g�~�P7L~6[��z�
�I@~�g"E�eA�����nΦ����U�S�!E~�+�"��ԖP�K7\��.��ڠ�N�DYoXg[FR�F.aȡ�0��ϛZ�+�����uUȼ���c�4���?@�H�F������IK�&E��]� ��;/�Z,�Yz�S�_���b�A�����A�4E0�|X����B��߮����I}r����C�`��WN.�wx︍��ٲJ��  �Ļ�5ؤ:za��XFO���l�3�����hXi�q�߬�.�-z�#���ݽ��t��4[��v��p��M@��YG��
?�R�aZ��]���ҍ���(bPDaBb�n���(׸�f�)�����rn��zz}3�=>��_�jA�n���� ��<�k��/Z���0��%Q	)�0�[����c������-���|5�*��e�Luy�Q����7q������E��m�J�Zw�/����iM��V���n��6|��U�����ڀZ�Bע�ҳ� ���rU��7�V�.w��_U/���j��jR[���=Ɇ�)d�Pm�����/*b�&� ����[����:qd˖�����`��<�2uTvu:��*�.�����yw��=G	��{����B��
`�)�P
A��_E3�w���M\ӫ�7WͿ�$̴8�>=��.�P�.����8���|s�N�;u
���1�K��N�.�3�݀��ܢi�A�n��t�iKp�Z^���r�ٵO����h�N`1ZC�!� i�(H�㗑|��5n,e}�=�c�dj(B�$ɠs�+��.϶��6����m�"D��mh@FR/�Sf>h6{X&�]-�~��l.�G�6��a��W����]n~�c_�_���%dh��H6;l��T��b�ۓ8
����Z�.�V�~�+4���%q����$rZ#B��xCw�{��<������:B�!�TqHk}�mu�Q�bV5)���2K�_�-��}{]���l�i!z�� [�RJ��cЭ�f��z���O�߽ez�����o�b���M��ܿ-�����(�lޛ�Z�}��8$kӿ
/i���=�ޱs6���L�8O��em~/��oW�3�)7ͧaK��w,�[��/�n��+�e'4��p87�Ҕ��)�&+��j�������4���<�6�_[o��~yۺ�\�;��;9r�6W�ihג�% ��T�h���F�x݁ iV�4��C�����b����dW>��4<��%h���k;�Is�-��������C��3�euZ��KG���W]2͎�Q��.�[��Z�:V_�Y]F~�5$�l��Fc�tu��M����SƓ��,ײ�&��������2U����q���0�o�.�m.�CO����*�ɺ�t�0_��oQ�����$�"Ġv�[}�
���2����ڐ����%�߯�@L4���)�gO/��Ϳ;�������R_�C����'߂�o��i� �LVpE�R��Zɓ{Y��V�~0�[7C��m}��FoR�b��[w������݇-��@}u�m&"�	��Up,�jf)�5Z(G����)!4�g�}�}��aO�H��N ��W�W�	�x��Ua�#2�Ԋ�~j3��/��WW��vϊT��dQ�C�^~�]�[1�Jh���YC��ڂ��M�~)�_j	s�n�SB5>���&�H���6+k<��)�E�Oşs�Ɏ���e��F[I�+�B�4������A���[�7�
us܂��/dT��b8*��Z;�y��Wu	����o+S����\�y2W�Rh��HA���W]	{�n${ݚ�
�=wc�V\�����ҷJn���|[�����B�;�e�υ�NR�JQ��|�ym'�Z�޶˸� ֵ�a�x���S:�b���J�[�o+RBeH��|[�y��:���J�kɧ"e������.�Q�襤��No<������z"G�N�#��[����+z8�BֲHP��s�Cu1���Չj#@�;��H�-~���f�_�]�&�-�dwVym9�RI��[�j�1`PC�X�:�]Ru]k��^�&?'v�/3�8��������s��O����wAm^P�r�6V�?��Z:M.�ۢ�(��({G!��O~����[�=��Q�.��sx5=N�Hl��W?�WW2��<śrt�����y�쉫�a�@�K2xAS-)��l�/O�j�#�`�"-� =�[h�(&d�B)\-g���j$B&BW���fIXډ}[=a��,�{UEt���1�j������t�b��O�p>J��c�G�+�ڤ:6^�M&",�D�Ǭ:����j��[��HY ��F�T�Ay&-2H�Q�͂�mל�|L#e���%�;���ڎ�>\F�||�<�U-3��u{h�b�����՗�;υL��p���ݻw�t�\�H_��)sw�#�]V��T����E��׃���ަx�7���h�"�]�K�/��┶ͽ��{����y�i\\�f��~'Ñ���Q���d�������|.1��@�.��{�fF���me.q��HK�s�!՞�r�cy�R�m�Qq���(=_���_�+�d45{>��g��}0`K%�mERh��k���,?����e���U{t�hP;��R��7�b����u�'�g��M��ѯ�<�t���
����K�%%�S+��n�s�y�a�'.��vt�ED
ՠ�Ve�؛Ou�C�c.T�]��Xz>�qn4�VS�G�a���L�=s�}zl�%��l��Ӡ�R^�|yb��{J=W��#��2�_2��>
s�z���G��i�ܧy�<�3��>]����:<��H�Q�1����z,�$O�@����ώ.�����@O���@���++��S���������\f�ܹ��������;��5�99���ܭù�.[���}����˘�%�}%��(`t@\6x��������"e(EI��&V���retB£��>����M���_1��f7nd��-`�z��aR�z�t�0]C�ȕmpG�c��+P���ϓJ��
��]�k�!=\v�S@�7���'M��;��6��\ӽ�w("+1��?��Ǎ|���3|v����j�e~e��y,:�6�rB9"����Ù��u����-��=����K�Q��<�5�so�^��!z� �Pjǅ���g]���@'&"H��E�g^�j�����^�3z�CN�������9�i���F�z�����QX�eG�9��4vw&R���w'�5E
Lw��@��'r{�ԩ1���3�gw�8;��N�!�_m�w'^�N.iE3$��3����t%N�.^���8�rpШ���n�|��y~$F������?��a�zW�pq����HiV�&���0��w�+"�Jz��7�`}e����XC�C��7���'��|��֧-��s+�W$K�����W���X��c(s,<�7h%�Nzb�z6�Qoc�X�!q�G&ǜ���r����@��i��7	�;�ޥz�x�|^#N�1~fff�d�����2FE!eT�ku���R�X8N[$�X{���ݩb�/�vƶ}W���>�&�E���}*�h#b�p�A)��>N0����f���nb��6�h�	��6Vp<3�,���f5橵���#��L�;0�����7
eզ�ԼNHt4��߃�}�+B������t��#���Ay��av�6;(�����o�����l5mp=QP���`ln���x���ڣ��?z��D��u�:@�pڈ������Ŋ��,��e8V(���]��Vz�\1q������pZ.A���v��~�F�[�.}NcmO"��sY��i���xt�-�\��dSs3:�s���U[��7����5��z���-��JPw��-�����=��
�*	��u<pB\�������qG�xa����r԰�יk�����.��((*�~fIII��=��U"Gc���@qsQ\uD�x���g*yҨ�"���un��e��O���D;X2���rq ��~X�1�%$Q\ڱH���ӹW��8�����6wt��E#gVW��e{^�C��U.q��:����Y��#�щ��������G�tG���x�/���}!��¨m�Hy��8pb�.���q9q�[$''�safe�kŶ��4����"�A��*r�M��9����C ��L\Ev\7��r�ȥ�#aH$�'ڢ3�彸�Ê4B�5��E�N��c'�!���xcH!�P�,&:1F��wG��yz]S=���;!�ӗr�I��u��t�ǋ|-�t�yz�{rr���D��jn9
}�6��7dfe����u�c&���58w�#es�Nb�w�+�;��A�b��Z����/�E#��<1h-���47�$�{��1�����o�\�@�̴��}��#Om������s`��0��V-K[0L�=���bMo�?���d�9ƞGE6o�َ�RM��V1M��o�ʜ0�qm�x?��6&�\�����<��K�iP��999� �ݼhd��Oy�]�q~��z�=�+��$������O{��/x��p�$ĥQ��svO���s��s<]&����U���3�V >�nq�5n��R���	���J����o����z=~�ƽQع�oT+զ�%n�@��=E�%(L����ʌ������MR�!��̉z�g-����Q�Fb����צ(��T�4�����yڟ�N��x�����W�r��\k�E��&�a/=[�u0���F��i�<�qI'�TD�$��^7ɣ��3ʰ�Cn�^��H%U�m:�$ "�|P����K���m�B-���Ť���{ٹ�/�����u����ւ�J��ٟq˫� ,�!Q��"��ث���0����\�C\nY����q�������C�"d�-�g;��!%%Ub��ۚ[�Q���Ǳ�'Γ�HV�ݎ.����o�8K��5F�L�y�;|جC&&M�;fܫ��ዮ�������Q���wm�&U�S���^����u��H<���ëG����rD>���j�1��}"���:�}��gƱp`I�a{p:!�)�$�e����Nf7�����1M��t�hg��9nv�&=mρ���b|���+H�f���S��|/����|4ʛ�v9�d�)&���
:��Y"c��44��dHgS]�&�Lے�#>J���ԛ�>X���C�(�Ԅ&�w��\�i��vu5�V�A�dn�vׄ㫔� �Ƕ�@'�/��"Y�Y^f'��
S�)D,ő�����piQ=(	� �����U���@�8��=9�����C,��V���B��@����eɳ���{
`�@����V��P��qt�*���LbUAg��(�~�ˑK�<B �����O��,����'EH�Ȕ:��`ϘOi�ɪgu= %��d�!1�����y���?#-�?ߩ-��9
,΍c��ov$Y>C��$��B�=���x��p̘X]t����X����H��H�\R4��q��mD�Zt�n��v�O��f�I"4A�P�%�\Rc���[���:
��o�q�]d���>��[���{G�/\�b0%yj9+�-R�g{0@�2�<4���j7�&`�v����!K���S���3�əB(���ǮF��\�8�n�%�?��B*yK͎��}K�i���br�������{�V���tؽ�Hr�+�$��4O�.`�-B����[���Ka��90�r���?����`��Q+�&���H��i���MJ�
��p����a�4U�8��IS_$�3SS��@7�ኒ;�,��q��s8���&��*�_�|\��.��LH���x�Ʀ�Av�<��;���o��
�z�g��N(K��[K2"I���sx�������(L5q>��1N�2��������N�F�`8aN��k�ȫ���q�u�L)c�X8�!�<�;,��#�uB�l����:�Z`qm�{���0��[q�{x�@�������>�����=X�ה{ٺM�2�PZ����<B\�Q� W��_��8���>�$�s7K�C���-�>}tp�蹻���FuBF��?d
{?<���e�� �r6[&���<�ۚB����ězk4���|Q��4z��+'���N��)�,�����H�I�sh�*HK�B�.s��[(��%,qkP	�<!���ɪ�0gǚ���9�u2�=���8+���y<��>�J!*��Bd'Kv��Hd_#��3d��d�"K��K
��$[Ȟ��d_g$;���Z�������y�?n/�ʼ�3�s�u]�:�����r�v&�l��H�ҙ�R� �h�	���k~��sLc��`T�ċ���X�x���	WӾk�8"fo�F�,���q�ϋ�--՝��ֳ 4D�VA�%IA,SS�:�&�|U^�m��P��8/9�����gk�sH��n�C34x�Ɉ�	}XP#?�|(o��D�t n
�M��ئr7�Phr�JӰ`�l�\�Ԥ���{Dp0�:��?B�P��f��}���E���i�׾�i�Z�͢Eh�=k�{�����I���#����'�7�3�sӉ��i��XW�:�>Cx��G<�<u��N����'���O��;G�}�K��8h�w�%D�pa�d�˩j��>�-=X ��_aT�"���U�]{�mU��%<�I)��\qɵ���M�>ʮ�8�)#}}2�.q����b���'��5fΆax�2����J�4��Zb��w4���{~	t��ԟY���B� 5H!�n����V�
FQ���<����A̔�*1(�Tos^�4�� ��I $=ӽZ�qm��gqX����\�ڨ�i�M[����=�0&H�q�1♛�m��P����Ǻ�/��^�\K���9[p�UHY��A�%E��'���w����̌��AϹ�1���`>�TFp��+�SA4�m_��ctY伭6���c�]/@��_ �=�"�����2搁���}��$ �G%9L�K�6�aX��)~N�b3)}E�(��M�!߱�R拢ܱ҅
�%
�v	�5ʠ�}nEGH�;����J�E���R����+�f 8tG�U��&��̚����~L(b�a�<~�C��~U���X�x.���T�/�?�	�izt���W�l�ͧ�5��˧�2c�#!�ǴG�0=��Q�lb��[�b������3��]�S\�d�D�J�M��lߏt2��e��S0%�8�|������RrPf����8B/
�d�gE?���3z��6:�W;���QTG>�d�;ՑY2F�Xg;@Aځ{�[��y<}���Ձ����a�d@��W��MEP����1����~���W���z'm��}G=�.5}_H9����T
)6���)����B&���uK��1<�wI#8�{��$P@�Q��o'	�瓡S�W�SW�w�F�p����}��ӭ[����:�e,�͆�4�4���k�����i�|��<��z�L"TSK��u}��N�O ��7p�mݯS����`�}P��cH�i�kR�?d�WG��'��3�9���n|hN�\y���|~f����z>Pl�$��� �?�s\aK٣^��� ـ���'4*�.{�p隨��6�A:;y;(+�#�w�nڏ�
SDj���a�`T�����z�"3�f<��۸�t&k!�����S'�k��<X�%VF'S3S���(�����\۹�*3��i��]&8z����P�@�̣q؉�L<����q���^�V0nOʨ!|��i!bٙ%;?�rt~���g働w��GEai/8$m��
��}LשN��ʞ� ����R���c�i���&jD���A�����s�?s���Q��@�?�o8�qXcBT�����d�����։�6�K)V�I5��t�#�&�ƌ8w���ñ�1��M�ڏ�G��Y�f�1����G�kW�+�F�$LQ�Z�ާ�<M^>ّR2#%� ���/(
4��Dc��3
�D��"Yy(/:�l �7��ue��j�=	Pr��b=�I}G91���
7�#;�������e+�6�
����)&D��+��l$���َ�)	E�'%M���-��������֎X��d*�O)�Q!����Z��J��[qR��^U>��&R?���z�{�cDm{㙈e�4a���B==q��M��13G�1��T�_�ѯ�j8^�P�B_%B�G���<����s=?\��{Q��a�r>���_����������Siu�)�A-m��e���~\X�6Ԃk�X��x��<Tr�.6��z�]qn�*)D��c}knr�d��3��l�Hp>>j�x@��=Fްe�AF��\�^� y�;�nrA�\��ǲZqJwB����c�]�K$���Є_����d���@�J~P�T�/��r�&�ّ�`e����%}��wB������Ӌ���,�"��*�?L�W�8�衬YƁ>s|~Ff�'�*�!9��㟚Kf�;�c�N���7�a�����v,>��Rxm.3�][��6:
��a���������_k����Lr&�o��S�H���v���߾7.��f%�扃������G�b5�[����GZ �ۂ;��;��jer�t�g�O�SeA��
G7n��V��`y�����v)�����m����O]�-z�b� >YK��M��]�C��?��1t'�����"���k�-�<u%{���5>�vS�hu��@¦N��<!����z��dN߰�k��P�a�F("l��!�������@��j~G7b'SQW�F��9-36
�87� p!c�<��ASdJ�!we�� Upjb�#�.Mp*.��Ԉ��.���{�z}�%���ׂ�a*e����m/`lP,�H�%A(Ǎ_�� ���{���Q�[�L^Z�6�B��8���@�8X��p���"gP�?�-Ͳ
�J�I�	��Z���'����D�����c�y8�kl�c䣣b��%?��DE�ϼq��ӏ���B���?{U�p�=u^[�B����:�QWQњģI��D�I!HϦ�ě�W�h@f�/�21��X���W���6J���r.w�A�7p`�Ǫ�N|���ѐ���bnA�}0��y��z��{��D���\_n�2c�gn[�+�@a(��z�}:*�W�T�^����P�{p��B��߰	����+��PY��ֶ2]4
D��A�/��G��ko�WIӞC��-ɂ'��g.ۼB�Zט��	5�2!���ČŇ ���Jz�8;X&E�7|;q����j>��
�3�R�P��e�	'QY�R� py�9"�>_s`�ü�E�?�NR�!�?��8(�$m�A����������*4ZR�м4!���"���������ӨR>�W]0��}e:j#�O��IK�`$��;���p2SII���S�$3�zu���dy8��a����Tİ�'��䂷ׂ?���|��H5\�\�/��hq y��i�fL荽�c�o�]j0_�:�]�6��Q���}��<7/m�^��
(��"��d+�/`��	-~E��e�Ӎ���,@����ۭ{�5��!È[���kјJ���B0��>		E��e��p2�ٗX�์��k���/�, r��*^�9tP�]�aN�V�A��~�!j��ۊ ;�9��ɣ2���M�
��Gq��}fJ2��nb�>����#�*��S��8�? ���Gu.����i������F�W?R��[����d���̜�\�!���b���l��Y8Q�9�+zY��b� �.��-��١e,�=i���Mrj��ynd��gqԿ��l�QI
�7:�׈ի�գmCeʘ��:"y(`%�JZ�����&5/�}��
xq�	=u�M��Ӵl؜ؼȿ�r�T�P��:�#�WkY$�.�� ��*�`�Y��n�$=$C�n)��CBϞ_B������H���Pd3F�dt)���Ӟ;?�apW��P��$O�yԑ;Q�WI��?�W��qDk�&�G��&K��Rau�C�)�ʔ���7����:��L*��� ��7�����_%K	��~!y��ډ�*�(J���$N�Y��\`���Lo�a^b�ÿ���&�|q�lLb�_2O��t�4/yђ�h��[�L����f��6���W�^�h�L}��zG��G�Ny- �ŋm-/؝i�
C�b/ʝ�����Ń�ec"H=�\�u8�妴{J>�~��J,n�F
�i�����O�꯼-w�B��E��5��>4sR��M��2$U�o���~�?�;q� ���@��!�]�g�̮�wҦܒ��& ��~���^H�#�7q�Eu�cp�Dj��w����t!.��W쭷ä�G����DA]���T�8�m�~��J���@�CN�>>EɅ�kY�Jkx_ �yq-��{q�aX��h����r.O����_[p�G������D�YO�7�h# ���.  i��Qg�'`���F���$:5rUBTv�*�4e婋��;A��߸�� ������"Ɍu�c��2���y����߼DҊ�?��߽e�E�D#%��3��(�`c$�>�2����>`����K_�{'�zը��`�<�4}R0Ǧ���oA��p*���ڴ  ?�L'����R���g��{/�^1bc@�`k�?���>�l 4[d��tM��#���7�X����]��E���gӅ
���U6�펇�1}>��I�6��?�D��`="��l����6���E )��eҩM��G*�/j���{v���5ӿ+����̽m�����i��NG�6i� :O�Z���ԁ�(�w�`[��#�9����m�W�9]��]RFjR�mȵ k�uyQ��G���Gi��.��e���z���7�)�j�5g'�n} 2&!R!�6Tkz�����)�ÏŶ��M/9A2:LPs��ND?�>�x�F�/�vp��g2G�c�,JN/����������R6@sT(L�}�2��Y�m}@���*�JG�~���޺u�]��{_�J����BUFy��4`������gFn�B=��x��Q,Fp����5v�Ӷ{�H;��������D�����,t�d�����s&cTk�w�#p�8���X�g�(�
o3��ޅ�1�cd�oԌ�}ER�{�k�ȉ� R��H���*��\|k���}����;�\��Sݒ����GX�}���I@���,"����)E5�C>ym�:�=��@)~����EKn�)%g�ݐj�y�T*���~�F����0p'ten�5�K޻�CI����-�J�8�V�=�a 3�`X�p<ٯ<�[;����?��^jJn�Hw�|?��e�UV �z� �X1��c�ӂU�&)���`�z�M�8�Ec
5Bn�T�i���'w$v����t�p7�c[2s�z4�8�� ( eWF{d���-\����y�!|t��{�D�$"��A�I�����i���ov@0���3����kR�D�)��B_g?�T�3~���&�d�s���3���e����M=�x9׽��KM"�&��Ee�//��;84�����`͟>=�`<R涐�H�Q�2E;��]��ET~v�ܣ)*�N�w�9��D'�]~� Q�H��Z �N�i�g��<F��`�
(��4͟���aZ��4`w�LOg���_���/��,�����z�0���7��0wT��>���(<oZ�RX)�y�E��� �����a/s�d�X��
�1�ޱ���'�g4��u�ҍkMo�ǣc#B�yـl�4��>�s�G�/X.�<.��i@ݏ36�>v�{ �P0Fٶ�wWN�O�x'�֎���i�l�s�@����n�:��K��)�U��ы=̝8�Ƭ�6W��p���tK�������U�{�G��q�\�qX8�?�H<��o��>A�@k�Xf�!�.�b�S�(DZ%�F��ķՈ�����F���dgw���vtsc�uY�-�bUљCue�f����LLL��h^6E��p𿭕�B�gqq�?���ٳ��� �c�����_-��7g{��� DX6fokz]���2�R{ %F�X�D��G4ݜ�H+y���[��V����mC���x(��:tI�혿&��������e��Jw��������y�FLV����H��@S=��_9��q��^Q�0��~�G+��&'BE��qx��z�%�
�9�Ƚ�#T� �x(=9�I�YJ'ÃȔ��TqVR�+*ZZZ��O���)��LFEH	�in���}!��u��)��`�\%yg<R���}��`oN8���_�Z��_����L�6�9�5��kS߸ʃOVV6�痘R�ơ/|��5�c�}�-���b����/C���N��� �C(()����+�畏�fU�~vF�_Ft˓O1�K�x5@ca���Dfȫ_-	ǥ�2
3U*!d�D��nY�F��lB��k��_���P9 [��hPa���p�ͭ�������A	25!�
��%c�T�i�r�t0��w�Y' �)��\O�M����Ho��F��S��n�iɗ�k���q@�+����O$y7OO�F��o��u�+���:B���__/o^:wnyyy����W����׾[=KH��U�0���˹nN������_���HM�$��&�w&�7Iz��tL�::�dx|�Hc���9�������vq $ ڹ�^vI��JV�z{̼��`Ӈ!�U��32.�dh
6߷��)Ѿ�t����N)�������bI�l$�p�S�����hy�$�s�:�)p�9��W�G,�,<�����kp��,�����!񻞾�c�ͳ����m��V���ܗ���MF?�joc�2ѷ��gt@��B���O��S:�԰@����bs���/�(`KqReK��0��X��7 YMb�'�q��ƛ�����Q�m�[DCC�̓�m�X[�/M�<7�ח�_�ݱ�C�k�0)�O�n�6�p�X�ל��Y(̧E`��t�-ܖe#"[����Ro`bCJ�z���e4s���m��N��q������F{���x�ץ��L<��|hmu�,!�%,�������Df��^�м�.��rE4��a���&T����(t@z6F��\C/�n߭"L<d�^��}E�U��ɍ�ME6-����g�aV-M6e (����B���{����*������"�D���r���P��{��s��2���
:e�.D��(�	6�6����7�#�?ҁh�A	s��l֮`C���y�z^?7Qօ�B����#���xU�$
w�>}:
������W7�֗�Y������Sy��aK@'.�ɳ����'���=5I�?[��4O���~�{(�a�����eSꇽ���,�e�Þ9��)�D"G!7��ń�� WL�)Sm�щ+(��o��������,|�o���+�v(߶5B����Uս��(j����I}}=��G3"���M�t�{��FD�WV�j�5�ͥ��3cDVIu�<s%����fr*'���iE��',����	=��"Rs:��֝>��^�/�GɅ�}�{��T�JA�E�}y����Uͤ* +�o3Ix��l�����>4����������c�R�es�`Jjr�����8ݸ�_7-c(���^j��KK���{���o��!�����Ok�,��NÄ떋��<qM��ј8�~�3g��ޕU��������(�;w�d���y�є��T�mX)���ϫ���	���ſ���%��UA���mwL��l�-�Λ��G�]:hӚ�<=�luP� 0�?�<�6檋���/ܪ������e�����' G<"^C� OAx�-h��[����$�^Zꙋ�� ��|:1`�^������V聞�G�ik��qO[ B 7�Lo�����@}s�z�Ĥ��\���F6ѧ��Cd��h�¡��9�鯓$-4�:i��iQ��e���� j����`'��"Oo���&��(M�\Y��W0���xF�r*4]P�m}G��:�U��������gn���{��]j��D����i�u`��%AH�Qؓ�l�"�s�
��n޼��S�]%U��U�����)���qJB �*.������Mt�J�d��0�C!��b�P:ޤ�P~����n䔪��܁���������I��<s_*���ً�����b<3?۳�^HMT�&ɻy�U��@��'R��9��Kb6���yx�?j+�?�Y�7�:���x%d>\�-�GLc�!�D���T�?~�X�������a"!n�2BBB� {�&y�����rw�7��ɸ�t�A	nB[&���gUn^�[��jC�zѡ��1������S�=����m�e([�����5-�gY��_�];��զ�1�����mH�Qq��0����o�T�Lb���,�Gq($�w·���6V��?��QD?p�R�o�Li"�	}��g�X䃃��I��£'@:��W>��?�8��e#qcx�ۗ�ʘ����h��W�:�U��\mU
m^��ilԡ����N��"k�x%�bu�W�ݘ�^G;tt@0�gl����QZ!��0����(de�ɸ}���:'c�оĈ;�J�,�����g�2$^?O:?��aX;�&%a���%�s�0_ȂD�TSp�Cm
�jB�vd5xѾ��9�m�)���Zu	b�#��a�KL���;�<����O�{���pp��´��2ﱘ��4�D�ʕ&,6�wf�ѳ��{:�����8���&A���Ysgx���h�p�p����,+�~�hű\���l��&K-_W	�`��/ޑq_��������+�Q��3Wݵ�!t�/�S=�/���$�XR�)D75]d`a�c�!�;B��ڊ8ұ�V���+������`8��xH05��J߉ �2(?p7�r5N�'�~�w��8���G��A<Sk��g��;��+�	˯{�c �}|�������??}����-��tww'�mԠ�w=��4����"z�(z��Z,�*�zd��_?x�nLAA�}H"�I�R^5���~�&��4g�̟���F�c�$%G�Zbl�%"��ܠQ�����u#:��y�$�S����覅>p@׾���κVz�Z�C<���f��;6,���)���G��C��3'�6� !�QS��^u��E
r�{ag>�]j�?��t����z�����x�ٔ�ο�����O�U�)555��~,��Z������A4 �R�!�݉��F1qq.UUU۲Wr�u/lG�aM��F4W�vO�~���[�����&dG�>95��w>%B����R���7������Ɠ��X688�uQ�ٰ�a�W�GW��j{.op����r�Oq��[��W[�+��(x�8uw��	��$�/� ��(m����E��P��"�1,N�P���|�Ԟk:EEV�t�ջb^M��$������k�A���]�?~�O$�hw�U?�7l��'�*�RT�}��}$��V0���������q�+���O�������X��-Yږ7n��<���?�T�ۏ8�W� 
�c�@D�$l�#��a��D� ���*	�mp����_
����ʠw( ��YQ#��;_������#�bZ��]BT�c�k#��`:aH#QFL-n�')�ܭ�,��j�� :�j���O����1����zI^ 6��v[kQ�p�w���!���-Ki����&�
��o�����/�������8p����/��a|���4��kW�yCF)�yx�4����1z�vN�_���J֝�aW�H9��X�� ����~��l6�=@aH��C���7�^�W�V����}��}�=�d���X[p
""��FQ�[I�uH��[���Z�s����eC�V�2�����#h�/�Uvl<J4�N%�x��O��
�a�(Pb7�E�SUt���eٿ��|!�\^S2�Z�@N��B,��)lRu#t������j��S]/�{� �A����K�?�F���������l��z���{���d:TS ��u:���}%uƶ�:��m�3�B�<���EXR��Ϛq�]R��%��_2)4������|Z�K�������34]~���eZ���Ѣ6�����B�j����f7C�_]�I\��Ѩ>4��*�o;y0�^M�V���hM"}�a��R����g�=�ZⓂ��Tym�yN����}$\�yr�o��R�[a�����᱂CA��\s蛢����3�4����%�9s��������I�C�@Y���I�L��	-�������ۃ�����o���'�"I8T-u�����=d*�f˰~>ߤ:��֠�~��
ύO2j!��г����X���|3Oi�;�K6�#���0����A�'����O777�E��>��/�<kMN'���)���ἒ���ʷe[�Ih.M���\9\p��=Q'��i�A;�	�dϪ�q)�+S��:ѧ�w�C�PD�WT8�իd�j:^̈́��Ukj$���_�W
~�6uA���u���#����	1m�O*~�fKJ?����AY����FVj�a3�(z^����e#pH���VG��K >�y4g��1W����3��g��FOh�#Դ�0ᇣ�������6�c ��7�t�b�J���\��c�j������8,�c�*���2X��0~���^��i��]
i��h�X3��q�7�����a]w�@�`jp�矕��^HyT4�J�@���'wҪFZpm�ןa6]����"�&�g��ա� �깸��o��f?����5��p���.��*��� ̻���T��6QI�$ �r���?�����_�|e����;��x�8iã*��{�X�4H b������������>-�Zo�p�j��7�PMMmt��:���!,����:?�(͘\>PlGn�<S?���Pz��� !��w}�GC �	�@Q�[2V�vZB�
�Ѿ��󊆈
� p2����AU͎��hL�W �5��e^FkB�@ߎ�uug����>����P��I1���L���5l��;������ڽaK������T�	��g���&�O�nf
҈������D����u�|������'���bRF�s��F�\�Ph@@�5����0Xh@�a³�շo�=Z�Ef�'���wP�v�Y5:
P�������-��2�o�e�y�X�_H��.V�'��Te"�<)�}�L�%�}4T�S�㍚�@��7�_ٽ!&�n�J���kH�˵x����q����o4,qv�TL^�h��
�eQ!���v�r�s����8~�E��@;<k,Y�^,�<Ԓ&��17�����=����h���{B��2s_��d��%_щ����V;g�3���}L�A��Ғ�Ҁ��Y*1}S=D��(()��ӭo&~��=2#O
w��ǔN��CW��,��
�m�f�|Q�I�C<�i��'��3�t���:Y1w�H �Gop6�A/3@�w�?���
�+�|���j^M�����4�>t�!�Js- I��6v����b�77=�ܮ�CC>�X|���������V�x���$x������t������x��]��C[)/U��;�v��
���ٳ�.�o�IJ�̖#�V�p����̠.TH.�ݼ,))iik�}���_Y���v2��'��'���m�n�2����@}e�����ݷ��+~�<��Pp�9��e&���z�kDx��	qq����-)%%��x��RO����z�����E�r��Cr��i~_�8���{h-y��e��62��%{���T���*ϗ1��$ v�EɆ�m���o��ӣ��cz��c�?z�ӌ2+b�ȑ#M���)��.���0�LR�;��A�Th����niiy�DV�j-]�����`B@�M�|��v"�)�O+~�j4�bjg��[h(�vѡ���~�%��"�0����J���W~�~�6�s�S3��a_�C'%��k��߽�S���˦�?�h�Υ�k��(�:��z�����{!����S-Fw�s�V(j�����Y洵�^�R��ީYm8^G>">1�����tY���(?����ux����.7hb����th�3 �o3_w5��6�;���=��5��R�.#�P�s\{�yNԀ�mᶹ�ʹ�&�,+4��|�vZES6Yq�N�����~K ^�B7Ҿ�T�qu|Je�;����uΖ��0��*@�6�Ҵ��S�OOFG-�����0��uqI�O�A�5����ʖ�����j	��אռ��e��BtѰ�FSLW�`T�5D%�?��"����7']�y~�,�?�#=��=M�2��9�^�re	`]�콊(ޫ����n��U59�r�M�ڋ�o�d���D"�</B�|�C�\@�DU�`�!g�-CI�·Ȝ�+�h/+�?���g��ek���,�JB���F{����}�$	J�G���>�Y�bG]��gP���coh��څp�wB�tɑm�!к�]�w_���s#��7�J����P�dL#��2~�L�e��|�[3C?7�Sv�^tm�O�QJu�r��Nj��n t�y+�S��D����9a�cx��8��-���c���A���<˯	��9υURJL'�9��MlY�wpp��9²X�%`/�P���lOpL|��2��<kJ	%Z��I�������M;�p����Θ��-�g��1�������(?�)�����̉�\�{i�Q6ِMț9�S��[���OB��|�F,���{���Ndo+��1C�>S���f�=`�(���{�X�c���<_Dm����=�b��>��߿b�S�m(l־w{r�|']9"�Kr�wE�ho���e��x�~Wq���l[/�۲�j��U��]A�1��̮�^���{˰<��;�5�Z7��r�F�)@�ƔgS!�qGn������A�Vr�w
�3r�xY�$r�pb%e����b}��ٜ�U�{l!Y���ࢳ��_��9KMe���!ǂ(uw!��*6p�'�FՆ��P[�}׏�%��S�]��H��ELb7Ng����x��@������E`�F"J���"$Z.�`gTioeo��i�_�QR
��	��vv9���H�{c��W�l���aԪ��8�6�/"��t݁�̅F2�����'B$�>c�x�%^�'���ZL_�f�\P;`r�v�->���p�\��sKA��@EcC���XF7�փ��V����b$�8/%J%و��j�-7�~k�UiԮ9ê�St�=�m'��G������
�
�d������%n�#�e�1�c����N���Pj���2��F�s��L�A�S���$J��o�m��mAe-�?{昁΋y�<���]?"�͋��ݥ�iX���
��k?ҭ�҂3��}(F�S�-T��szUG�9��	��9�}B��PW<T� ��N%pLjz-��J:0��1���ҲJK~�>�eQ�t��زP��?���˅4~��u �[P�1������dl��X`g����W�H��3*���$Kb!�ư�t���'[�nød*Mc��j��*���q �M�U�i�W��8�W�_k��n������z,�Z�jO/ia=�W�C�����"+wg�g%������T
�g��W�Y2cM��:cj=��>�YGbc�.�888���d���*�u�N�k��k�޳�MGqfU���_M
�fJ��?���'��+�q-ɰFHm���9�i�L}b��������~��Z/�h��8���W�,z�$<��PS)P[[��<c���_f��NX������N���5�*4(^�ɋ;� �Bz�syUp�v>#��U�]�.��=���U��e1Ry���1�Z1����ku��k�q|:�+j��J⁕�tړ��Φ	��������ޝٞ
G��Z\���{�뼪�3h�	H{��`���������'��g� x���뷝��E������z�O���\���i��������ʖ�c�p���ȩLNXa�~v6J�EEs��B�Fم7Ż�n���Gu������LNfJ�ZX��a=~�nm�8uY;���S�7�S����"����I�����Ĕ�L
�aTT�����K	5�u������$/�7<&�47ݼ�L���L���Sw%&�T�U���k�?�R�LXXا��:ط��N�=]�u�pT?;ߤ��<����C#�N`;��bA�ԔL��c�$H�*��qX㣀�Ä��@I��H"U��]hn&��j=�.ɟ�	�����P�������j����v6��2j��9j��di�ٙ5wt�q��X�D��(��)��i�����a�h��?w�6���vиybݰop0fi�e")��}Zavvv_

��� #	آ̢RaE�"�0����a-H��g?�Ι��Sv>Ր�|������{XZpa�B�35�4PC;�f���!��:�}�}��큽���4X�1��yL�Y�3��3�1��n�'^�.����!����Տw���J&6?�m����;���iW4���Q����P#G��l�X���Й�-'舄M���ភ����bbbZ��~l��u-ϒo�_�<�X_�{_LKGgem�~��r�,l�t���=ő#��Ҍ���yR���l-L�ìy$?����U�}o�9恖[6o����|�M�y�$���������g���XO��.l�\����W_���-�9���_>���r��c�X� �K<h�I �< p'��l����������gȼ6�x������~o8�uc�a�/
�rr����&g�t���/՛�P3l��kI�S�<)�����#��;��N�2�'EZ�]�L˼�*�R	�~
�q������lגWH��_���`����L��6��XA��5P�;�x�pL��C;}~��R�Gul����&΂����VT��
Kظ��z�@@��2QyyA&�=c#�ԡ�p�j�b� ���������J?U��dS�kmr�g��F/:-f����RH%��h�۝M-e>)�!��\�(w����H���I������AQ�4���[������[[Urn�ONc��4l�Smm��N9M��E���_��?A�K�R��2�nV<P[gQ�x��eA�?��l���FX�"!!Q��p����zZ�8\�
�����p�������G�+�t�X[�?o��Ÿ׻צ��p�����\��T���p�e��b-O�5別����a[azP���,�V�sk�~�f����Ǭ�^�K�`ȏ�zG�7�Z�wݽ�gH&�G�_~�'iI�������W��a'4��7~���^�9��kD�������XX:L8�Wn�ވÑ�*_�i�YX\t�J*x<��rs3�g�?���y�������r�[X>����z�<��m��^z36!!��P4#�<$Aj3uR�� @�p�5JU�s�㰂���rS_����_��\9c@䵯7#�1���J�D���q.�gy �������;��P']�I=�{y�*/--m�׭l�{K53�Vw����_(�l��GJu���Ns�mjB%(��g��x�\vɚ�����z�#��C��~���8�Kk���W���v&Nt3�HIH,��Ok�9��>���9�d��4�U>d���,x<>��As��C�$x��(�%b4������K�kS��[���vh�)<!^rrX�����c{�"���Y��P-�WQ\	Y�Ox��zho(��1�q�N���$� '4�e��}���H�B�y.��	.�8��֖y���+�]w�^��/"g��aa( ��8c���!#=��ފh��B���%�Lug�}���,�������"�w�֓W����5U���}zX��1�ݖ�u��ύOL�5^xR ���d���!�}��?���O�@xc���%c�_á�#߾9^��܎�������v�H)^
rJ�ߣ�(xݫod�dce��8�s��ʣ��l�Λb�1��brr�7��B��U/�P�!�'Ц| t��X�!�����f�+{*�)Tx�Ǉ�FT�'��C�^�����0aD(y�uy�V�ަ��z���7eAV_&#�/o��-Z��7Hg2��p�mо�D�jâ�8��F��}%��"�%�'Q�a�#��a�%	�v<�����5C� �	j9L�Y5<�}� ���.a�js��4C��+`4�}����^!AA�F!�n��'ON��T� �:��vz:�Ǐ�v��3�z�kj���T�,�, ���I�<��^�xzg��#io2P	<g�c�>B���ZPo�ቹRM'@@?c�^P��k��!n�vck��,]�6of������8�!�K�Բ���ne��乂��<Њ�B���}&8��POg����xi�5��(�@��ʿ�;����U �ą�1�0�TDAd�pH�?V@,֯-LPmVߝwH��Ҡ���������iK����S��c{1��1�I�?76uui=�@	�c��v�kk��m~�|�B�����{�����/5������	�/�5�ӁKKOlJU>�iP0T��?�|@����#NBsuO�m�L�j��1ZCC�c��^� t��<X���D2�5������ L�{�:I!����͍+�b��N�rW�clB��-��0!�6ˢ45�;~�L��*b�.��B��&�IX�I"�e=��y42��0=6YA���շ���0kY3��L�m�rT�m��A�JtH޵�_P��?���2p�0݇���r�ߒgbҐ�t�
���M�㷳��Ru��<"@Z}_W��C{{�o+ǎR�@v!�q^Ue,��^����tOa���Jѩ�~P��׈�ZBJ��r���T����r�NsS�Qc�}�?���KR�p.t��tg�����cQ��=Q�$����I
�������լ��o>G�#�d�Ör��ʟ�!n���9����H9�z��g��������
�2��SQ��zЮ^'8��DN'�(NZ��?[G�a%��9�ulM�MR�8��Ng-]���������MQ�٢F}_�<�L�U�gqq�,�O��у^3S�s4��6�����<Ug}���n�����kb����%�� ��ٳ��99???��@i�|3��* p�:�O��Bsq (,]\���5ή�zB&U��s�
��sl߂v$�?VY�]ar^��W-R#�u�-�-zbf�E����̓�僒��=�α���#''��P�(���mX���r��x+�9��[�����z��D[x�G	-��ж�yA�/��{����&Y�)�_F 5��ۿj����(�R��6�n�-T�T[:%��\��9��x��.�'z:�!S ���c����n�|o�4����޾=�����zq��ΠZ��QE%��w�Ew�8�_��/x޸����EɬLG��g׶�N-
�ѹ��FD�>��B�4��&NC�x��1#�å�y5��>����&�tX:D'���m_�Z	� =��q����Z���b��קWd�g� ���x�YPW��0�ȋ��n%�u�"�O�c��V��+G�k��e�K�Bм� �5~���0��E��~n�T�B��;�]Hh���O��L<�N�Uh�LV��� ���f`k2uM5��;F�_�Q�����B|���Gٯ����Zzm��L�>E�����w��rKCN- �?�~n�X�5��t�7����(;��в��N�Q� ;o�3gz�猾gF���;�%$8��l6mj*�O���"�`����Z�)��r��u�URv�$��Tk��}@���a}� ��X2��C�Mg�8��)	YRR2
"��B�b8������׈W_��B�Y
*��3zB��$�뺱���8Ol�=(.��Q8��)�L�ƾN\����vϻ*y���5KQj��ǵ!ߵE�\?r�X8U�?������U � ���َ_��
�yh��W���q�*i�}39��a��D�S�'��࿳[߾�2��2������~	�������Q��}�#ע���r@�s�%�d��\�g�%�x���+Q���H��r�\���{=�8��!w�$^m�������c��H���q;���^��7���g��a��s���[[���Z���XRR��8�baa!�'6��-A�b�[�w����  �q_�L�ό���S��R�2���h�.5�/q�J��	WS=����Q�� !�~#	j�>^7W5"4����39�e��r�c�O;����mma���������x�6�΂a�F�s
�d5����?�����P3˝i�}}h�l�˕��8LX�-ȏ��j��+��v�����uL��),�[�d]�oLu��f �ra<�H_P�i�g������ *�З�o}f��Z�¾: ��{U�2`��D��� IEr$g�)i�K��%G��n�Q�A�w�A��l|����8����<Ϲ�9��LÏcc���8<��m��힛�{P=�"�Ц9�K�{��M�p_�^6o�|,�5�K�����]zx!W���z��>�7jn����E�X�&/..���B�*�f�fhΡ�5ax����AAuS�7EZ����x�G^���e��������D B�j'���K�h�h�9A�,�Z��ma&'v�ߦEy=���J=���K�D�DO��V#�F�,_��s�- ��[�l,���)�O��n������nU�wHu1�� i�j�wx!x�󆛛�.��31��1����z=&��!A�_V=��� �J�[���߇���0�(הmA�.(������윴� @�/����A��o��D���`ove��O	�Pe���5!���P��e��je���C3�	i��a��o�ɡ���֎��.�`o�$�Ms�W�y�C[���,�c�ݫ�ɻroj����g,�F��k��e&Ӝ������mN�������9�~L�*�K%�K�]�������Jo�;|qS����П<�����9��r�g�� �ċ=e^�d�:ku+a�߿��������>�0`U�***\n?�5���z���|���%��v��:�
��K���N�N�q���8P:���/Qd�j���Y՜� ,�\�p�8�X�0���xs�.�8����+�.k(��e��DX��ݍ��R�R�O��8#���.4���`�YL"�Z�m�^���`U����L�D�7�)�k^~��9��g�����58��s�AN�©�탐Q�{C��8���o�_�~�pprҁ6g�甖s�Tj�4�lH	|bO� 2�ϲy<�@3r���~j?���|��999~n�n���}iҹ��墬��b�5�C�Lo���wk�V\ӍH�/��E�V����$��w�*����Kz��A�����m��,%�0Q�B�;:h<�s<����T\�TT����w>��L�ϗ@k�~��꫻���I]]r���n�P55z�iW���;{*�X�k^?�����t���%��W��p~��n&h� i|�d6m��i6�{
絊�N )Ay�⊏��UJ��oe��šn=�ͳ���!�Kv���(Q�G99�o���',���=���%}�73i��?;��PM�Y���w��G�TCz^�O����mӑ>K���ne��¼(�o�%k���j�̥a8_L�=m�+3X0袤z��Y89�,l��i�������o i~��&�c��SZ?y���?+W��� ��2�����r�-��t��3O\�8ΆǛ�`�R�3��':, 2����V���J�W���RQ�Z�4Q��F��{�������1�k�{0z6��Z��"���Zڜ�����_�\>9)hyU��f��9���PP$#:$�o��\�ξ:L/���Fڳ.�7�YXY��A7�7���c=���3i�@����޽��+AC����cpN������e��~w���:�H�U��W��)�p���X�7;�|*S����ihhlBD#�K���l��ڱ	!A�i�����*)�� ��%P�R:.!���7��m ����pl��b�U-�[,av��(��ju1��ѻ�/C��t�<�#��ǩ�uF����{*fhre|<�ҫ��jz������
e� ��?���:�����P���u���ĺ�:K�%���^'��o�%9#e/�_]~B4W�}�n<�8)R�EY�n��K��.�T�^��s���t1u~5�8��i�4r��{��݉���kᔔ��;���e9B�t��.p9b��lEp;j��!�9�U���o�zUY��c�	`6bO��GG��G`k.�����?{g�/� ���<��"����w����8���?�:UJ�k�[�pz
��o�&��x	j�J;�v��^c���Lh>�s��ׯ�m5����>��/�M,-�0��#�G��_Jȏ����þ���4�׉���g�="9�!o�rCc�ߴ�9��v�.dZ�l"�l% 9��xi��H���7��Ď D��2]v6a�NP���W��8]�*��F�.�@�ր �j
:�D �
 ��*�J��'�_ K�J��<@�������Ɉ�IM9�������aa��m�Ǘ�0�[�oj"����6�C��&�p򱈡ȋ7�U��ݾ��H����>!�K���)YB}§N����G�b0A^^fp|�  C�_=:53�7HctttY`��mll43�}x3�U#.I�řt�t�`$�ũ��q'L�T�*u��("�O�F������<�[����o.��P�{��}[־�A�>�}��쐴ۣ�@�@h��x;�E�iYQ%/�	T��C�������ԑnV_���`�-��'(��A7!� ����q23Z�S��i��w�/S��^Cu�$�
�����r��h�srr��2�mEZ�Nݼ?:$j��>(�,���M�ڕ?F�C��5=�|ɇh�fk�[�zI ɧ�eg������`��^�1/��>g(s/2r��̻s�ʟ}�K��Tn�X���S�7�r�Y�G-��c9r�6M3En�ܷ�e�r$3q��~|��86�_R� >D�S0�f5,�3�}N�Y��q�m�%�q�SNw�;�M�g��ڱM7��^�tm(��yǦD�M~���&���k�C�**In1B��ݻ��3���i�P����̡*�W��ot��5ǢGߍ$핹�w߱����}��.黸�p�Pu_���R�ڡ������'����[�/9����0ş�2C�?��򠁲����ڪ���>k�	<�m���4��J :����E%����s�1������>���!��VΓ�C��tɧm]�%<���m�$N��'BǇ�#�6�����W::��1�����x���c�΋~#[ �s�c��lll��s���v?hC7!�f`��T5��u�F|NjO���{�'�X�>��N�̧�'a#��&����)��}$Rα[���ﻧS��%%(�EK�*�>Y[󵴳{r��&EeC�����a����:�Hy�2����`K���t��Z��ݗ
<��_p7F�nd;^@��y�CZj���<_��"�g>��>=Q�U2~�^���Q�3�Et<��0}M����9aed/"^Ӌ�����keeUYU���???��P�#�w|�a?#*����ϟ�LN�S
��<���($��x���}��3ֵ�9U�ɬV�*`��͉n�7Q�wg�pt�DS\l.L>�ڪ��{�2B�??��l�+ϻK��4+�\bD�$�ۗ`�D�sr�^\.�*T���v
~�v�3X2FFF�7f
��	�p�>�k�wzZ�adB��D:Àtq��選D�]6L�5	ɦ��ak�Ⱦ�A�A7kz�2t	&[�������pT�lA`��aҗ��uBl�M0���E`�^\���>拱Y��g
|9���p�u껙�oK�5O��X�x2��EѴR�R�*��j�W�%�}�5��K�Ea⦚�],���(��@I�pQ��ɐ
sCJ�s���(���~+qZ���Mh_��cS�C�za��P���w����˴oX����~�t����UK�wݵ�u�"�R��2��wml<'%*�����	V�R��P@�ѲzZx�[��!���1*�I�*/�a�ᦣЭ��#"rғ��Ź�Ѡ�=�hP"'z3ڞ��=v7�/+Ҵo(`4����Zoz�Q$���T���aDl��g�XO�����,�Ͷ/���x�$�O���SC��Q����o�
����>h��*4��u�U�/]Bl[89��O��1md�OJ���3m�;X7�=
_�7p��v�m�Y��..�����3O����/�&J�2��`��
:A�;BP�С����GO��b�}�H��7�2���C_-�¨�z�R��w�y5Y|�����i�0�,hn6o~����hW�v4l�|�5�E�����s�>w6B�i�������0?��+�b���aXt�8Q���+Q0_�sVgW���=fi93܄Tm>�d�$�j`��&�-z��,1^�E����� �tu�5��h��>��kC"1�<��0��H:�_Pv
��o�S'ѧ���?�����4e�|Q��R�u:�`F�Xr�5
r&c�i ��Db��M� X�O�۰�ڳY�4��6J��v,�2?�H���}�\	�@����9�\���8::k2i�*DG$}�m@d�?��BU�DNe�Da��d!��M<an=w|�O�뢇�=�͉�o%���8�ΔQL���a'�ƹ�E?n�@�T�oĝϝvB�"�����NYt�!lt�y���Li=xBq���Dq�prR�;��S|�~��X�2��{��	
%��T�%�����Z�������ށ�n�%jh$�hf�!if��=Lz��R�ϭ$�FϘZ܍6��٘�Z�m{��/Igg�;� <��{�k�íҏ��^�	�_�'D��:y��`]��Ȁ�~����)a=Zg(��ɑ	&����R�T����
�3��cF�\��>h̼�C�;<��,!Y�4,t.C�]��"���C9=299)��l���NƓh���Ц��]�&	�)s�2vNל��I�-"�ͩJI��~L�y�'6��(~&������0Ty�62<U�Q��58u�ɬ�{G��3�<��<�p�4�Z��c���'�%�7���"8��X�A��45���2�ǋ�
�D��vOXp��fO��o��t���a(�E'��v��0Ɗ�n�Y����@�uS�4	���̮3Lo���ڇ�'ٛºҴ��	�ʡu�=��G~��M7_���-vNľ�����fS���w��[�8�\�)�z/�AOe?�Δ'
��1��j�'L-���
����`��6��DJ�v�������~z�=��["�/�x��߭O$��շy�����mu~s�.�6*�ah�o��HXj-�иu�������@f�F����g2��|U��~�_hb<��ц%Z2��M�͜�X:Hw�5��b�g@�ㄪ�᧚���e���瘬�1P|�"w���j�Ƈ�d�0��ペ�8�Z\�*dk[ZJB�Fɸ(3���V��>�4$0�H�t̔�-o�e��iצ��8� ix����HZ:�Gm�ո�����Db��L����]FwsBc���Y�]'��`��#��9M=8%�������Q�)`�^��HN��t�`���/"1by'�S�U�7���3�K�Ҹ;t�P~{��b��!�/b
��4)QS�'��<�~,�m:�(�	q����2�����h�� ��;'5��ŏ��w�����y�=mGA&�< � Y�)Q�-�E��/7�']s��t!��Mi_�;�W��.�(^9=��`��q����%<aVŉ�RUE������e�A<�_����0�S<�ܴ����!�lz��A*�m��i$g�3B5��'	�f��s؜֊ej�[@>�c{~2����n��g���9�;���\��:�9)���N�uM���q%�?��x���,_�):���IO��"����Ԝ
�� 9�,J�f�8�C@�CQ���n��^|�r�<��Co�긯�倽V4���A�Jx�4'�Y*�X(����[�ƶ�5���c��[_��)F�'��3��F��kS�ф2�-��~	_㕦=ՔD{�'�3��uV��������3m�I��P(��m��C��'�V�[�����W~X�ϱ̳�큚p�?�J�T�h�'��x���p���!��R�z��:/�,���B��#�(�v)�;LM97��k��K�ڕ {'�
��DS,6��`�ԫ���e�x�N���^��+��X���#3��V��<�l��	�֮�	��kz�6dZl�J)�V�d�61����I�؋����s��	�������<Ut�4�in�\��#&���?ќ,W�!�����Qs[���q<M\/�y.i�j����6t��_{F�Pyj��&�C���r<����.?�_0�������(9f�
�]�����,߬TCBB�k�U�w��H���c#��H"|��� �_󃕧��>�o���	f˫gc��Mz�e�r� ��z	{��K�t��P��08�h[؛��6k�a�LCI�8�t�s�m��|�r����v�����c�hǛ7�������{!�_�#���O�\iap��j�Mc )�1�A��+?gP��N��	�F�1��#7&�WJ�z����~�=֞ ,�ڵ�����])L�m2��"0�U�q�k�ٹ�HZ����w�X��v���\VN��ƫ�`ee���b���[fR�o��׶���l:n|.���A��r���EY¥�5ȑ���b��Wy���+#�!b俈%%��8����ӌ��>}����[�|vכ
���4���L �D'OPG�,]����C'�b$l�������XCF�(�p$�($��r�cdb�n���[7.���t���d��w�*W��%����Y�s0�r���	4 ����Z��[�u���;�>���Z�������lb�����V�~m���;I�.I��h��Y���d���K��N4w���H��Г��$��|��/w�(�hr�]�|�<�Z�&O�)g�JJ�SS���Z�I��X�/�֕I�`c;V�b0��ASI�ɕ��Z���O�xp� ��J��/J�L�#�b9u��%��qh�* i�ќ����(�ۊN �c[���bh�5����n}��889���=���+-*�R�]�������x�2a-����Z�gϞ��?�E��e�Җߔ}X�*��N��;�tp��Z:o���j�q���?�@tq���,Z{�j�5\�0���z�-5�lN��X��t^~m�B+  ���Cl�5�+�÷�`�w[�$�s���T鱱��,}8l��C��F��@�-O��/��͛��=������)T��v����4wt���7�q��b��-��rz
R���HHJ,<S���Y�[@M�^"Q4;;�F<S��
��6q�b��<`��&�2�̔r�
�~`�""Di5�D�_��"J�}�bᶲ<��H�^�iO{�ʃ�XO�)�56���6x$EIT�)q�,�wj��9闺�������1l��`���ڡ^E�6�9v��/��wYZZ���j��L����V%�V��3����j'�7~��as�������F�PLu�iM9����E�^&."�jßY�T���wE�`O>lU��u�G���B��X��
���`'6���zҟ/sk����|�FD5
�����!�hs����{����qF�(�k?�xf�����?�y��x�,����Ϭ�2Խ�ԅV����WL�
ǭ�>�H��nK>��0v3ڙ�h'<��I��G[[���G�˃��j����[�kq�<'�s���kqS_O�U���cp�q����{�f�;�u�J�Ȕ�s��sނ;�.�/��/����S���	>"`����m��^��d>�w�^�62�9����[���4����U�8���C��J��Z�9@J�Qz�=��M��ue�}�T�q��P%�X'�/j�%�-�/�z5�@J̮������������՚;���n��)B��k��;cߍ��(���'�5��5F�r�ҞM ��%q}zy��� y��H ��xN��x�Q��A��~#��{�p�?�PM̠K�|��^^]]]�F�9rGX��B�����������|>�*Z��1D�dP�x#�K3�Z��D�ߠh��P���'O�ެ��ߵP��T�k�?��?B�u.S���O2 '���g^��Ｂ+˿��.x7c�>H�ζ��2b�6<��a��PVY�In��#8�V37h�����H��$,���im�jΒ+�`��)���4���h�f؉
X�k��E�f K_��iU���t�-��Q���E���+_z��~~:�9����01��F�����R�+1}


��.���c��nl����N��BP�Y
 H5L4�{�y�6kTE��Σ��=Q��_,��{z[s^�ܱKCw�S�C�"���:P����lg�]�J1޿2��|�V��֔��^[@#��%�-n%����Ǌ��Te��P��:�����D�1�-P�l�"��c%�]�Rn�~����ח���$���,i�&һ�:�(׎/*�Fw!}�^�U�	u��+�2�/� ��?�@ޤڧ��Rź�9�������wQ��Дs��>���xи����c�L��4gL���/�T���^&�6�;��ǐ��5���Gt��2�l�ۻJ��X��u��C�+*�� H��)�I��s
	ɭߜ�� ��{/�i���c���b���UI�tK5�,���?����Ӛ�\��c`.�;�<�4���8��FY��n����
^�o��x��s�׿L4_�ǜH$қ�Z{�ͿZ�\X����V�g�jFm$
����b��_�w)e�S'���ȩ�ڕ?N� ��`lxt\Na���> 2�'����Sq*��'`{�<�<�p�~���)��0�O�ZZ����,����%�"�����`q&.yz�2q:{��L�j�	*�K�l˯��8g6��&��J��t�Q�"�{��,��ꁲ�[�:���6h'�.)����eaJ�p~�yh�i#��V���ՄǼS�o�e�I2��Z�{�=K`y���������_\>u!��;ᚨAVc�=������kq��Po�ϒ��E'ȞZ�H��J����9�kFO8/.��N���1a�����u���/��Z�^v�q,���S�� �o/�5�S�	�*u>�4鎸��{*i��P��5e���yp���<�������V�5��N����e�{��i�X� ��$78fW�܉�(
�{�0�_��ѿ�����&TDV�
�퉛�2Tr^@=���E�%�M����<���pW�=kq�,�o�l��N�ń��9ԽQ�<�͑�VWt�Aب��x�Rx��C�t9�ʊ	�e�|��$s��W�,�Au��v�	a�8g% ��F�
�LT��烿��'$\��ǧ���Q���@��{n%�{Ny{e���i_�wf�ˣ-�	�#=|7V�������(ܮ�w���l �Z�W\\�  ��^�fc��C'B���n4|ͦ������\Ξj(���V��?þ�?]�����#��@��'�ji��u��'��:�-��MK�	\=�Bu��D��yx��j>(��_���b�/�'ț�}�ƺh��f��s=��g�;�yd�Pfx	#�9\P8H�w�����g��k;���)4�ߢ46��7CO>���H���cp���`�U��&utNgy8�%���r����w�	���$�F�� �1�������\@j���Ea��0�.�!{[B"�1&�@)�	�*Lc�h���!#���-�A������.�u�O ��Ӻ�����h����F���oE��ܾ�$��� �u׊.+:%p�'�����s�ǽؚ�-�ʦ�T8�o����U�-{��{D<5��Ff��
��Z���i����pJ�H:�P]�)��-�-[��k�;;;M�,om���b�E'GG�
���v�b�)���*�:D�c�m�z֣� �[�@63�5۾������=ذ'�����*���Y���$��_��Tg�s��Z�"���jQ�����:��9�g�����~��[��cKk��V͌��'�J�kc<U�j��5�����@1�(1�����5	_#������ĩȖ�WWSs��Vo]@C�s��n� �m��6���%V$��@7�jz��#��F"`Mw�a�	��E��.��rQi�_iI�I�Aa8�&�ɵ�:��/_v|�aZ�ǮA�
�"ȀaY����?��ʌړϙ���0?�nv�%�АK)0<��Ȉ��[����Y�,OP�D�&�ZH����#dt�G]B�}��G�F�-J 	�nL�⳴yD̏A�5{įc:�e�6�$����uuu�T�{���A��G�6]3^�࣯u���Y"�@b�X��0�Lc��=~����(�lSd��<�1�=��p%�U�L���
�Lk�0TŇ��fБ�6��?�*�?�7:�iu�w��ۙs/^��a�%3*
�t6��M�SP�����΢����g$2->>�_d�_���Q�9yh�&��ԑP,=S4A��{wd�|��@>^��a_�	j%��|��/m�hS�R`5�3b�D�{�����Ђ��Ǌ��5F�i�@u��H�ў�C���"���j6g�\�l����nn=mm�}�9 Ո�<zE!(
(E�r� �5K��2�,N���MM|K�晬�:Gk����{�A�-��9�ΈHvU�#��R�R�RMN���
uZY>�D���$ݍw/M�{��sru�u�yS�:=�/�&�W�Sz��@p-:�g��֏�v��#��v�kmm��nr��'>&�����En�H�U��u�?5rŗ���Jn|����O릞�O����!3�bN1!\I�:Gg���˽������x�(v�:����d<zĲs�ࢌ��#C��;�P���9:�S¢a\�Xd��c{"������[2��AO��pv\-�X�ݜ�?<?�#eP�~Ùyma��ꋐW i��8:y�:�x��3z"����H�����WU�h᳧����6���!�{�÷j���kp�Z�R�Ҟݝ��[!;l�mQ�������G����9�22�o��T[�H^�A��(���#IQ���'�'����i i13�ն��"�y�z�?X8�d�?VV���4�WN1Ʈn����Ƃw��8�1�]7�iۦ��nl[�^��'󢬬8��P�<�ng0s ���o���LD�U�n8�e�>����Ҍ��k��H��tK��������Z(t�"�ëk�?����E8��w���g�F;�[���1fcc���6��9vCݲ������ϼU��~랣���Q[�l�Q����)rF�i�u�܃'H�J ІŋӢ��1����&	��Ky+��ñ�m��%��z���I'PMZ��_��I>/+�k��{�����a3uKy��=Ւ��駘l�L �<%u�0���lR��/����W)?�[�'�����$�%J�����$A���P1�D�̭�|���2~`fe���p��/(�$Q?�(D�Ȃ�ޛ�l��}���P�H���̣��9��$K#�"UG0q�Ew�
Uqs31�4R]�S?��4)�^�{�ZX^�uu5S�W�r� �g�e,Sgq�Of,Puk̈(�BS�/ �]­�Bh�������vf�,�]���T$��s�������c�$Z�����)�=|h]2�)�g�gd�u�ţ�����&���A�z� ����rU�Q�Y4�>+��86����\�ݒt�A2j�2��p��Q�F�ie�V���KH��0��* fO�F�p*N�5=�(J��2�J]6Tyx$U�[g���.?��F�� ��_Z��C���ɟ���d(�� y��|W���sOǉ�踟����Ol|-���DMU �A�f���N�o"�΢����R���$�t�L;::z�������������42		�U<r̐�������.>���T��N�6;��~�J��F���*s���8ȩ���4r�P\l9ݷ��#H|�Q��@8�	Q��tr69���~@�����m�ݵ����I9��0v�a��jd����D�����#j�(:�13�5��]i��;'��1�{���V�]�L M�~�d�T�� hO�L\��#T-Rα�s�=�ޏ����,$'3g
 >ϭe���ޥ8����Q%�h��.���,�a#���6'�)7v�ʤ3�UO��|�&��������
�����J��L�����&��-�5e�Cu ���q�9��N} �;{�1�D<����e��S�?T��*Xk�x��%��k������å=&�6?����>bد���W_!Gj�"1l�k�'a7������C�p��_�$J��BU1�$�撗����!}m�*VMŻ��e�|���Uܙ�3Ƒ�?��2�D���k�[�ng����p�D���z���&�_gse�~�ƒ}T@�ص����-�O�^=�Pǽ���c9<g�y��0A�=���	�?��,%���� ��Ã�,/#��nAL�߭�(	s��A����I9҃;���$c��RL���N�r�6�.v�<�$Y��T�5�Bh�	�A�}�W-~��4)Xd���$��zs��f-.��a����21o��h�_le&���tb������֌_`�۷ZW �6m�b�u�}E\��8���5�o��Mf�=���Ex�S��������O��vD�M�4��q���S�MR�1�0F._��[���=T5]>|�@vnnE+�f�I^���i��$��Ȯs����g<FHU�,~��'�>T}�S�
:�&�(�$$,�=��϶����VM�	&&�����[��b5��@�Z_lE���	�齭~����P�Ŀ.�wi	���sv��RZ�u�F��;Z8(�����D3���3s���F<ܞFF���ж�<��EM��������3��IO����ҏ�<?��Z4����*��Yf�L�M���2#ߋ�"bA�]GXǆ��9�A0hiUr$��*����B���ۺw��gK�������.��n��/������P={ʉ��4�>d㏳��o��	W��q�Uɳ�-�[DG�ys��C��Tf:ۛ�8z��Vl��>���VVD�Suy�{�U�j�E~��c�o^5ւ�Y�-��3'ߔbm������
�*��~��O�����S�t�z�3�_�H��*�ɉ���0ɔ���������bi@G^���uЎ��<�ǌ2.��9�_�Rk�_�r�æ1b��o�_s��Te��CC��69�x��q�jA������"b��2d� 틱q��Ϟk ҷh���R��T)�	���i���XQ��_�V�k���C\e��ժ��g`�`�m�j16M��@(=J:���:	O�|--u��'X�dp~��)R��bO���Z����*���_3d���,�"�'#=u�i���a�p�˴X�|q�2�oO%�桢*ыP�W(�^�*:�r�d�P��bf�E��/�3Nf�Vyf��ks?�u��c��I&8�������My��e^΁���ɦ����
d�"
O�;���vBx��/�'u��&oЍ<�1qY���w𪞛�XhS)6$�0��~�?�)|��F:[��"�¹�Ƴ�TZ65,�r>��Y ����������(�W#�����	�!�;�p/Q��;&+��>�1)�l��c���G�!�z���MZ���M�X�>�)v�u5�v�������[&����Y�I}���k<E��"�Я��9�N�����D�z~���5�8�̥ƚbB�'!�ű/�k{yٳU�h�)���b]��O<5�tP��3�l��_�	�vd�epgO����3oC������W�T-��-by��=���'��d"Ȟal�Ȑ�҂ٱ���^|<��jY�'���4��j"��TShx-�ie&u�F�D�<@�c���1��Դ�h�Hn�Ɛs�y��d������߰�1��0�	�{��E�wf@�Ǵ����mw�ExK7O�G~I�j\�J�ф��<S*�:A*1E�dM��zv�(��w��5�h{���r��͍)�b � �>bU,�N�.��D�u�p�Dnp̚�w�,Z�C�d�Gc�r���&�W�*����0���<�}�S'����=�x�ʷ�\qjcZ�1�T�6M�
��;x�ɸ�JB�6�¯r$u�_ˑc	��?��
��)R���a�姗�T�6�膇���)��]"�"Ӷ3DW�M�]��q��ϴi�:�}5]�i��CC�73pG�6e$�����,��]�a!+�.`��]��972��s����R"�h �O��\~����~U�V�L�?+�E�1e�)�/o�
��Nn��Ko��tL?�Ms�B2&[�D�L�ev� �]:v����ZHԎ%q���a����J�6����=�^�����4�^z�Q��HڃG�xH���IoJ�Q���H;.��������؈������F��*�/z0��[�~9�����v�Κ2|��Y��Y��xW᜛�Y��&�~B�js�#`c�,g� y�ܸy��@��l����r�RT�R��2�J7�?-����J8�l�U�jY7=G׋�^^^T:.���x��S�gDD�
�ݛ���V�s<�8��TrzZ��Po_\ۢς����^M;��m��-/ 1��$�R�m�z��	i ��r���/�?�?eV��1p����+�)��--���W���c��!���a��䳍������Y��#s;�sg{���Cq���IsV<�/!9�T�(1��PC�.D?!"Xܫ�v�d�hp�>bq���@%
����n�u�qv�|��D�썯�xxk�a����r3A�������P�n���4"\;˪~.��U��%-���Vn�3+�T�
����ޚg���qU�ڤC�Y�QlꝟN{�3��Af[��j�������e���,R�׷1�¦p��_,ʺy��볔坞&�6tg$��. "�c�2�e��訵'�<77�G�6W����S���Ƣ�4�|Wlg�u�I�� =��!G�+vs�gE㓗��j�����<L��z�m�@�X���'
�ӏ9@E����?�zb-<<���A�:�Q�zgε�!��3���V�z��i�����#�y�n"D�3B���dq���pY����?q+�9�TCJ
=��|vF&u2�Xǯ���o#.�Z�%���4D*��C��$�=�T@���jq"�{���4ɑ��w��v*s'�_>�i$NYovd����������Z�}���Z��i�7��X/TF����W�R�g�����jZ��Xx�E��@��g�D���#�5�{��;;;\����"?�Xx����ҏn�1���0���yr�eb[�䜸�������4�c�y�QǇ����OƼ]<��1HƂT>_k���
�L���XEC�q�m��`2��7s�����(�1�ǒs��p�,d��[ngJ#�����e�9������Q�-?�\5�0 �(�X���J����3ĩ�F�};��:�ZT�OE������	�6k�>q�R	�Ӟ�w���t�^�	�+yt+�%��v|^��پ�I��mY��;����C]<kXe)���c�]�)���/�N�FWT�ga�
���'R�	�[VJg�L&����U�}�C"'Z`MH�^.�}m9�z�/fH�\���/̫#,�=���{��N��A+n�?pM�w3G��-���`��usV6������auՁ�e�n��l���-���gi����OTsK�Ip6iT<[��W:��/)P��s|�8m;c����}�b�mz��֒�ȃ�����<K73I�������3��SF&&��bwȕ�ݾ�U��G�ޚw�>q�8�⏫���A���ׂ��[���g�H��"i�>�\�|�X�vr�A�_V{��Ë���u~˼�Y�[��Ė���A�ۺ�J��Yrj_�upJՋ�2�r���b(�0�/������1�I��e��`Û7o�������nH���K�2e�U
r��	�[ �sCۥ}�♔�0�#/dJj�d����#!��)T<.=�3�N%����mz�{o^���|{�Pt�C�}����ٚ����=�����3N>��8���k�܇��|N��E�8���-P-L ��@ꗼ�a>��;$�~�9��5s����2lB��R��������ǪxlqͿ��Fߴ�(���/J��}l�Kn�G~u��~��VEm���M<��c����	.�p�6�'}��:����Ć�9i�%�s��7%xj�i��nM:�|u��1�����W?v��v��.t�o>  �<�a�#�"ߎj������?�LЙ���c��>�y(��j����NC�G<|�D�d��M�ŉK߼q�i�&씕�$����������R�������M����}�k��G	yy��'��J�g�etL�򻒨�K����A��Λ�CP�c�U�,\8���d�,��z�~���O/@������,�W��W��,_�+7�P>b4|�uPj�x��rk��ˏ����W͝9��l�M�j�˼C���(���	f�z�z!z?�M�Y����E�Y?O�*dS�} ��UՐr�a�(���^�y3$$���_��Qr����+���[_-��O�T����w�/��h\/6Ѥ� ���D&z�}p���Kc�W��LN�E��m/�g�������hgX������o�C����

��,�~Mw	��{g�l({���U�Ϭ�O�K6�2�x�e ���/\-�ٵ9��(�Ej�0���u��#@o,^����5|�J#�z���hn�
Ď[�� ?�/Oa�v��&�?|xx)��7ռ �ր�� }DVȆ�ޑ�"uu��]O�ꝡ���������.�c�"}�i����yV���tڻ'oo�K�O��dnϤٕؾ�C��%�]1(4��a֖��k�v�ז�����b�	��E���[�^C�К]`ʡ�;�6dT�u��T���Y�L�����
2�j.��p�_&ԇq��`�)$�a8ngWI1h;5G1ࡈ�p`uuu�œ7����}��g�Y�i����'�N�o�<��R��2u�Awww���/��������o!���0�L�~��������N6�%��^I����ם��*�O��Ae#�
���N��$A0��t��?����f��R2Mp�����<��웶���:�{N���\�]�ۤwg�� �&$$,(�:�����"�K �ƒ�xo��|R4��K��q:j���1�l+��w(���awjq��0LA�FL��?�N�ZO1�:t{��Z�@�!-��X�v�<����	\@'H|a��`��saBl+o��v���������]�עR;x�IM%��F�LH�eLc���������~�](�1�xÚ����mS\1�ۦ�i�s
$�i�U��l�[�{e�N����!O�j�䎙+����Eǆߌ{��V.�	��y[v����}~g:��sV���E�=m
o}8debά8�R�#�����׫�:3ޯ��s��E��0���0Yȃnee�3ו���s���J�O.\Z�r�􌎎0ق@�����[�B�xи�>��&�?5���,�n��8�y�h�#��Q_���������z��Yåo������������!��u՗�$�zW�1�[A��F|�[J^Bb��T��06���M���vcw��n����ܧ���.GS�L�����pM�2��q���>&���΃9��Lm�������LP�'����O�ux��q	<!pYi���2���VV�����]��H��媙���

��ӊ� Y��D�k�
�{ ?�����ώz88����E=�E�j'��P9%��N�u5#�j�JJ9��A�a�Ʃ ����Ɍ�ӾX;���x�n'���ή��'��zb��7�m�r�؈���P���2�F�����e���d_~�	�?dgs�H�^�d{7s����]��r=Q ��/x�hD����?���?0<��?~��_����/o�M5��/�*q�_[㭁��Nڙ`�����*M�:|���0��(���[XQX�����.��k��?¾;���������ބ��ޫ��H�BqrΑU�#+�̌�2R88I��V�q�W:G��~��Pw���������q�=���z>_�y���3��R�	�����n݊��떗�.�d6g���L(��2�����F,�B^ ��ۅI��2X���XfyKO�rTu��MΖe
����'�(=�z���r)y��n/�K�<Z�ey_�|)wd�� bg?/��u�YXd&${v���%M:l�}�M�64t��j��}c���p�&x�e��e��b���O����u:S+���&$����s���'A�0��v��X�g�?�M�E#�c���ߘJ|����p�����|�iVS�KKK�s�J��(<����@=-5�����)��o��7Z�_�V�zwC%���5���(ڠ�4�H|�0�b�d)�~=�圔��39{��嘚=��Q󘔦�K�/dm~����j-,|����*ܜ�����$Xgf
,�l~$��d��dȩ��k��ի�
���KK����]��	'�-�7�}ʪ�)bG��?{	�J��Oh���W�f�du81��Q1g���p�L'?g>�K.�u�B�z�5��>7+��XQPճ�&n5��I��7MOB��H�L9�-6~�O�H��W�+�i l��H��'��O.Շ���N��x�v���
-�b(;x��]�&�*�h
s��͋{A�O�0�� ��T���q;�������ԁh6pdA��ϭ��`޼�=B�(��S�b���
hDu����d�wT	zOM�^k�|�ا`S�`�ɝ�XW &`hq��KϛEe~�oP��&v�����9w�\s�$�:�;Z��w󌙀� i%�'7���������.G�-��!1`#���F���Buh�X�ֿA�Q<hQ��d͇�F4�N-mD���Q��P��W��
�5J�u����r�,����j����lm��s4Uش���b��ha縏%�fa|�M����;Ws���VW���e ���Z웈
ET����<��TG2k�6n*^5N����>�7�i\�/�{��z6[[�V]X��"��9�:ׯ¶��A�Y����0A)�.)D)���������aVN��,���fy(�hl����ȜC�N	|�4��k rV���wă�������յ5�%��J�⢒� 	����U��)j\���:�I��p��+p��e8#]VR6v&����x^Fg�7��λ�������J��A�e^�%qS�ٛ�hX�6K�����'+G�Vb�ԜJO�xW���Q
��j��iw꜇����Z�Q&���7|�Q����Pu�p�p|���|���d��bmEl,�,]�LNR��p��Pb����2���6�<�|v�'�R��?:9,�E��� ;i�NWp$�<E�m� C�j�`�͍"��e�@�P���m}ENV1f��\;�K����׼�\)?����+�6���r;s���lp���K�t��@���p0�D��H>����b'?��E�W,eDqx2�OMkQOT�<yru�k�8�N��*������ƔI��{x� �,�/N|���$���&x�Z#�d� ���1H�k���-7�"w?p��Z9X�K�L[FT�Β��OZ^����� ���M�t�\���k5��@�Ag 4>M�z���mR���4.j���i�����J�����Z���%���[q�G8$k2�!��0tR���a��/�?�S�� ��v&\0�K:}Ë}��D�5
P�8�!&_F�W�շ�k�$��ܜ/���a7�/a<}-l�猡�n����A�^��	NyY��R�ٸS�:�� g��:�Q�&O�..m(�U��A�詐V�z!ƍ���{���3+ա�����w��(� P��?�3�r)IĨ���ÕFx�'�yV
7�&KA���'����������<= ��j��٬;�Rq���wx��^D(w�=��X�i`��j��E�PE�	F����T-	t�<��{�U�@c�a�t0�N�����w���ֿݳy���A�sk�8����K�c���)�c<�W�#��k��Zx�<�>6֎�$�����+0�����rF)n֋�����L�̣�����m���v)���˨�*��l1��Fa�֨����xҾ����Z��h�"# ��� q08;f�sG����t6<!��--���?�4^9�N��^�/�Y#ಱ�[���}��PsGo��&��D���t �Ǉ5|�F+łf{�����jr�YV�>&��tT'E?My�N 	U{�}]��Jy&�������/	0	��r���]�۴@Hr&/{��3�KSD�v�)�
1�7�y*���h!/��Q��l9���L������}��8�3ښ�ժ��:�.D�[����q٧^T'�wY��pk :�v�J�QgtUr���3�\����'� XkS�}3���C�bT�21q8�e'� r��JL^-�:u`5���# �z`,F	�y\����a[�H=e��+��⻮Vb[k(�zK�<"��� lXe���A�f�)�0���Z1s���>`7^��p��-�tr�If
@E]���<���n-�|��ؗ	��:� ��}�0^���l���� W���o�z���^"t@��9߼	�� �I�u�6�& `���S��쪰��{��3a�y�����J1)|	���77'����O���C���Ͻ��\�#�mMǡ�\�����Ygw��G���g�aL'tf�_����v��{��'s].�����5��@Aٚ`��L.�����5�N��u��a�73����;:���?�e��?��:��ఱ!�t��sDs���C��9++�'�w�?z4<�����\}�(£}��m��Y�C7��W�����7hܵ��e����,��7(#+�lA��O���J��r�Qu}�&�X���z�.��>�d��=s"Q�+�:"���W���a6&f}�T�2߳<<چ�nfW�ޙ�$�V8�ܼ*��r��e/���ɒ�Ok�Ù�(?�@�� =�~�s��I� ��'Z�wz��m��9�a8
bxL�r��{E))��[$��+��xX�N�q[4�3[��]���W:�VEmM��y�t�*�M7�AxG_��à
z�z��(���㷂�Lkp0����S�e�ܲ|\�؏:�o���/�$�Ō�*a]Ѵm���	%����8���#C���m�N���=�<+�h�q|��o�*eX�4T����[]�q�u��$>����q����	'^�a��&�P��h>���R)��A&2�*���ՙ �r��
>�loػ�}SI��p�"�����`504F���6"u�؞�E��<�RG��7$��[�(��Ø���Q��/_N��EV$d}����6�D�e[�����5�GVOi2�U�I�"�R�d����D@��u���'|뒌��
�u[�%�����@�:�VZ����s��g�o���t�I���7���
�p�,zT�;qW��r"AOJU��,� ��2�I�r?� ZC�r�ꌟ�����_7�4��A~��0D8A�dϙ���B�ˣg̔�]�L�B���=�'�?��=�8}�4��o�a�&Л_V�Y�ܐb5-,��bR;��ցL�L��իWR�c\R����o�-Jī��;l��K��Zi�cE��&��E*s1J���Y��̊R�B�Fb���VO	��*��A��_
��]y�����h�*� 2��Z1�[��@c�~�UC��N�Pwl ��G��(i1�ժ*����&ܦ��c8���g�U%�$bD���*��n@4[nq�(K�`�mf:K�z�ٽ�<�1s�	zSɚ>��F.`p����V��@hb�
��&���~\�
b��WR���/
1�:_j�cR�]�.�Skz���������a��i��]ֲG���B+-�*�@$���_ �BB
��:"�$�s��Ta�Hs<]�}UTMư�,ؒ-�.J��,uGo��U�SD�}�GS�F���rܖ��
-�|r	�X~fo�%�Q&��Xy�KY��?Pwr#��i5QB �}�$y@n=������t��C7��>�G�!�ԯ���$�s�A���`�ݺ9g C�|hh�����,��K�M��r����ڟ=I(�e�f3�������ؠ�I�F�mV5ֵ1NH@Om���׳�_�K��q���5<T��2V��V�N3��\p��F�U0�sz|c�ls�r�<��Y�u����A�?+e�ʔIZ�Tlǆ�� �8_2�P�Sze�T�#�\�#}K�>��o�O���+�>��ר�K
y楙I��e��I�wJ���������%��=`���)qZg��Jt
ʾ*��;3JG��7���P����P��|N.ÿ�����
͍d2��k���rŝ��������,�KnJ<Lw��~V#�B�)��V,t�1缍�~5�xT��s���_�ۈ�'��T��f��yO����#��]���4��[E��?�t���lr�׉�ԃR���_D�$�]��Zi������yA>�8|N��OSS�Bm��A�.1� �iV�	{�ny�NF��+���pJ��8�����9�K: nt���c|R���Q@�����H��5��r���c@���	�]�r��<�F;��"���Ý�ϩ�:������0��*,��;��k~����\&+�~"�~�uMd6��{��Uҫ��|�q�����k�I��y'z����ԝ��^�l���0)og�����_M�l��9��+�w�1h,R>TL���?�q� Z:������t/�O���&���I�o�����:�Q�L�Cƕj�[��C��	�,��B-�����nL!�=���=Ӆ:I�`!;��r�� -ԧ��"���o;���gĦ�\��e�b`�4���q��kӇ���h2�_�u������i/�:��,��q8��ic�Ӱ�&�׶?�Ak'S�'���8��� ��>�)��a۳����V�u����+�y��łB�@�9�D��]�Q  ��q�`����VI��Y%	:9�9Mh�c�6M	�U$��J���#vV��Nz(Æ���M�E<��,�f�K�����Ԥ�XqCe�P{nxx�̹��~����X\,*f H�Y��}��ӣ������Zk.���'s����
�8�n�:��Oc��?����I f_NU�q��27_��6�Qa�T�{ ���/J�Tr
��(a�{Љ�[��%a�~)���E�I����(E�����K����S`�u#�<Ņ���]��M:�t�TJc�L�� 8͈u%"@7IA�q����R𯉧�$�+
چk�.�8L���Oņ�p��;�?�6��4�裞�h���*uim��MQ��Ӆ����
���m��㊹Y�1�uX�^Y�vK��ʐ+�4�*$��`�����
P������3y�*�8bm��I���*x>5��8	�|ȸ�����׺g[�l��ܞ�ɶ�X�������ё#��V���	��Ր8�����k~����oKԿ������kƧ��i4�v�ֳ2u;|�c?���I�3�b��{�����N�_�B ��y$Z7����N��_?T�z��aĤ�e�||Wa?�Ac���s�3sh���٢BM&~q�u���c9��,z�TA��=)�3}���용~��Ǻ�i��������2dO��?`?�N�w7Tl�>X8�7��ǐ�F��CF|���v94ri�D��=�Im�?S�P&�r�/��j��;Ǚˍ5��4����;�b˧�<6\+ �U)!�����܃�G� +�I�T�B6� x��n��}�q�E�DH� |ӡ�Y�PA=�s)��8\��#�J�q�j�z�ld�ZJ]�Sش��5m�I��w�i�˶��4,��^�'���<�x4��M�Z�O�+ա<2<,�hX�gS�Zy����_�m�
8���ę\@�U2��Ku�8��w�Ѧ'�L��K���t��^��z�F�z���ˈQ`����N@15I���ߏ���{��+�q�/���Yp�7��?���@�`�?n��g"1i^�|2�#����M츖��q����7&竬�Ь�4��;2�#�[����?G�B oh	x+u����9�nǱ�cB9JNz���;;�����,�è��DQ�Az���ivAĜ,kT���X�3===�D���&�S��3rT{��6��ݔ��(y��a���#�h���|��{Lʺx�o��6����]}�܃�����{���EgW��&�b���(I�b("��cv|��{j�	������`�]�:�mO$����%� k^����Qss������^�qh�eoZM�L'&���'�M�j�[����WV~���~C&������$%��D����NNN��@r�(׃T6��^�ؒ�=�ׄG�GF����]�Du���^puoytx�̹_3����|x>�[:n��ڴ $� j@@ 4vվ��9S����9$�P�2ݹT`�.�Qb�3P���	4�:�ƿ���[i�u���%"�������ׄ���)�8� O�9y8��Q��Ɓ���{q�=r����o&^Bo/���"s�N#т��\�����~�鵝�/),��M�6lX|ۛ�ɄF퍸(�L����@���c�n
K.��H��Q�h�7~�0���}��Q11�+W㘋ĵiw�V�zd	׆.���2KQ99ȞSAE%�[T
��N�����]�P��(�e�}��e����Ґj��U��1�z����A
���u8͜�R���	���?����Ȩ��n?dT��}�i\��_k�4�V\L����PQIɅ�S��C��c@��w�)ٻ������w�x��_���Sk�B�9�� n96�w��PLXP����қ
���*IO<L��' Ūqb�5�RsA(���fZ.�e����\>�GQQ�2ͮ+t��ьkzxa���z�8�{�����A��:h�,��4 HjW��`�>���`S��B�����Ҽ���a�ci�g��à<���ze�J9^'�
��A�''fW�ز��*�\�Zo��mn5K@��(�/A[��ڭ���>� �u�h�C�g
(�=��=P ���Cg`�s�q����{���U�T<8�W���^��J>>)�.]:�t����G@����z�ŵ��b?(����T�ؠ���69�@�bz7���M��/�έ�B����#�7
�Q�T����24Z���r����5�)��|N��YtbC 5����NL�L�f�JnС�Jp���A��O�D�v������-�N\oT܍����s�95-�w�%f�5R����u薦����$vg��^�vq`�bx�m,t3Wu&,J)�O��c,�S��{�u����G��_�e_$��r��Ǖ��V��XѷF������v�׶�й2WK��W2�> �M��/�������8Gh����P�İx\_㯁��fӭ�D�]������^���!�ڡ䄝?S�p�p�	&���������O';�{{;�;G�����J��hZ�����8!.�Ш����R�n75<n���
����D��])5y{B/����r��F������'
0]�����b�����Hu[rI^��LtI�!-�a�Ӏ��%��%�kǾ�ӰB�?q�|�㹞W�N� "�`�����*
Q��T�_cL�c��$2DS�S�.�JJ9yF&�>�sh�r:��Ĥ��U�z
��>�P��Z���4q�ؾ�;$X�[�t�Q�ؐ���/����A@wK���J,Ҟ��kk�f��HBEs���i���p]Ԗ�B�Q�;;�H*�ځ�A$�� =L���`����3��2��L��]��5G�g�Ol�v��LGӊ�ΚD�;�lV����?J�F����:vvT�gT��Wd�u'��f�~��P��9~���E4�v�K���'��I��r�.���~q3+|B<��7�$�lCq�S�;�[~ދ�5>kb����6�t���l�a�5��;[��<� ����c�x�b��m��3�(��tcWY��%GK|��<CT�C0��k�/0����e�	�{=�l�(�/�P%�zdsc&�>��&?�A�*�	�t�����l�>T:�sX�|:F�/P@M�[��|p��dk���B0�?V���}����?�<:pbv;O���^*,�ѣ�y�YKKK�?/z�������&�+!�H�d��� A�>�+�)��n��s/���46���p5�ۯ��1�Uc�ͮ����
�nv�h�GUתz���S�_�Ʀ�c����p�$/�X%�{�f��z���+ [�/�5�pW-ѓT��4�� ��9[��
Cx���x<m�}�F��YXka��]}>�����@ r���;�A쯸3w�ˍ'LT|V����������XY�;�� p3�$5��U��]�h������/d���,\�^�	�l�n9�`㋑�����m|{�>��E7�z�|�,�fa���ڝ���.3$�8��!��7��} �uV�Ӧ��G]؆j����({S����n- >��?��,;��ٞI������鋆,FXz���N��F�i���	`�c0mV��S�[�����8wy8�Se	ܪ��X�zvGٞ�JN����36K��ş>�(�K�1�(/�-���Y��g���h���	�eک�Ƈ?����후��N$SM�N�n?|�*۷����d�Vd�-kp)�X�K��LVюi��¿>y�XI����&��d��^G�I��i 7��[�]�s=Z#Sm����^�=�d*���2�{F�jU��/c��g�ȚwM$2I����Ȃ�y��1U����a�2r/���o���6r���ZT�4
3қ��wo�`�pWK9�	ǩ��p \�WN���XL�B��%�?��*6"4�՟��x&��i��~F����0�A�W�v�8oѯ5Gm����"9��Jes�0�{�eȵ�:xN��"�s��/�N���]S��!?Ӗ�\�C�-C��^�rGS�)HKO3�VH�~������}���;L��;����7��_�z�����UGGm�
���vmm��ꈱT�������Hq��&�ʒ���8|��ԼWpp}��몮6u����7b�&�.�j �+G�z2U�$Ymm��7��xv�Ȗe_��("Y��4k�������~����>��Ej��� ��U�'U��5hM�)���-�;:>�K�'�m��o}������M����˗_�z��as��7�KF��o%�w����G�9n�ާ��V��l��Tz�T�}�A{ZZ;�3^���pS8fH�H=y��'�^�3&5�`�*Uf�Djp:X<l
�YGWp���^9vO�loE�;M�Iu<|������@DT����>3�KbA�$o���3ޡc{ew
���S���ss���ᇀ�OnE}X�������#��{�� �}<x�a�r�Iˣ<u�M���`�>�Hi?0bY��o� ��I���q���>ŭ�ă�!�e᳹`�;�]M�vqumC���T}6�7�1�<��o-�>}\/E�����a�%<7/�n���8�cc)Tu�yY^~�����<���/kj8���r����x�H�a.��!l@�n�f��w���لW�[/�d+O��=�}>�Q׈X�r|%9)G�dn�3�ޝ���CO��ff�|�M���,�& N���MM]��Y-LU���-��B����;q�喡��8������ J�C�S��5�¥��ü+]Y��0)\a����l�dm��`\����\��Q�v����kJ����>|~� o{�+q�v�����
��p��o�`ű~��~3��P���H<�����ʧ��v��ׯ��W>\�����V��B�����4���8k����z�����J�g�5�0L��Vb�ظa"�� ��K4=o�?�H��Qռ� wE�]��-��H��9�@�Բ,��j�4r�ҐS����]�����<}*��c����bNEE%�*��q����ǳD��ځr��u���I����r�r��Q����4���2f��R9@�.z�|�͝�`+=*z�8���]YQ%m*�;�b���oE�|9�k%V������E���w;;�H�+ɲB�C�Շ��@�*M��p��c�A��7��+Kv1W�׽�;��c�#�ڭ[F���;�7���OuvT�҇�����K�A���$D�-�]Q�Bi�����->Ț�&�zK�-V�%K�L�V���uJY9M!��IU*%s�Ť1���]��7}ǃ+�k. �p��~N�6ԏf\lSc�Q}~r��6���<?$mak�h{g��J<�'�u�P�\�qy�/��r���fG#�`O��=tbqxF(���`�ނj۩gY9J��ʏ���4?�gg�hqf<Wҡ.6[���X���˱��{��Z��t��}�ǥsss�]�X�6x��r!|��ʗd�&��>��F����H%�e�����#�[E?VJ�\���7��w�`��`/@�1m�
����ex~����~��O7E�K��G��q��{��sRȠ|Ȇq��Ȋ;u+15�C��N~�!�6�;K?�t���v�R���U��j�&usA͖���,�)������H�Ё��QQGn/��Y��=��
�u�3�2��u�ǿ*��(�,�&��}�47�9���p�ٱ9�a�#�V8�Ny蟓/��'5�L���[�7�����1=}=�!�Lߍr�"�f�G�/^1�O~��63==Y��9�vg���˗���$��:�������|�O����3	$���`(����ҝ'-���,[�XPz.��#o����w>l&��8;�C�ٞ�a��7��5�ڑ��Ԝ������U���*-p���و
}��ѣ�x#���M��ׯ�hqn���Kem��tn3��p��V�;��P����Xy ��%@-��TF��#��@3)*��������'�U���G��7:�j�0�؈V��[����zY]}2(a߹?e�s����Y�e 8��l�i�r�amy�&���N"s�HG��@&6TD6<dbS�������W�(	���[v&�9��0��!>�GC6�!7;(��O��`�B��^�Y��c:�b7�i�b�n��P��X����r�*)~^
����?����B�q֯��qcT�(�Y�١�E�cA2!bd܌�ؙ��a�W�qš���s`�v����(�b�)�A�����b�j�����H&�a|ѥs*;�U���RU�93W.,�����7n��>�>�u����zr�.�p��
k�@�����3�(�́�Jq��"��Jga����|b�����$����YwC���iQ�����X��F���۪ۨC�
��-/_�V��-Z���é�x>)�&��J>�&������7`o딻R��[K��]pf���d5���gG�*��[9A�1��|�^�|�:��ϐ�(db�WJ�s�iQ�����L�a�' #����*N�+K�Q7��[���v������9����c:�#�B,��p6�D���� T_���_ُj�͂ �|~&>�<'3|/$���L�q9\�/@P��~
������~r�QwG���¸$������,�Ǿ�pMY�s�]��� ˌ�����[��;Of��}����q"�u�)x[J��' �Rvt��?�+�C�bN�������xB���kŻӕ#<*,E7f�c����}]�T�0�Ԣ�SaV5=<�껳1��~�S�Y8%d;�� KP�8�}��%�]�J,˪.�4���a+7���u#��mșԋ�0�l!���T�G�]�)���	CC�_d#�� {�+�DP�W/@x�3��l�Q����Dxj"F�ѥ�����ޜ��f�?a5I�g^!-
����$��з70,`m�FX%=������L��jnh�(�J���υ��	$2�%V�da�_�<k/O�6�9��򩑻��-�3L{��|;oq�E�cEM��F7[��`1g�����ʻs�N6B(T�eO�)�c��>{��a, s���x98�Y'�[<���E�������~�lWMĞ?���\��#�y7f��lRVJX�8����S�K	E���)L��^R8ߵ0�u��Jc��q�
6T�D�O�0�pFXtJ/7�����7 wg�h:�!���K���6��߽{�Zt`���w� "�fc����������EU��O�<W\���1��.k��Մt��iZ3u�5\@�0�r�>���-+�5�
�T�u	�$������J�n>���<}����Ƒ���tK퍝{�N�mssηg�P��3Z��QTTL؉���.��oe��u>�}U,���뭽�1�C�� ;�ʈ0<}�ݻ��z��%��ѡ��7oެ�gJUD�YUJ,��cRY����h����V �F?8���땞{�*W,�w�I�!-�3�%�gR����60kyd��ڞ����%a7ً��P�� �n��j;�c�������	��BrW�"�Ó��b�mA4_Q8�a�p >dm�'/2J4�l���1�!3�����i6���t:V+�[8�P䒮�Գ{ �^��T6z���{$i��d橜�W�xפ�­�=tҺG4� �y���w����ܶ�K�G��i�ܵ3<�ďf0�f=u����8{)
��+�؀˸�q��|}=iHB���q��J�OME��2��=7+1���kj�C��kF��o�O$:cWW+ ���Q�@4�9%b@c�s��?�����޸J��i/,V��B����_���=�,�י3ݵb�����-O�w}Hd�Bc薀�_pR��(���҈�hj:#�"����& Ez�J��mB�[�:�}b�D�U��Z������ړ��=�o_̅�p�~�B'�U����5�<�0��܀-]����7��#J�}�#��:+�d��B�U��Ƃ�36����W��܇
�>K��i����:� �����H8xŷ�И��ޮ�t�Q�{��]G=�p4�>�ّ���T���]p�0�1Nw��9W*ks�8$f�YZZ�m,}�qk0���`�G�K	Nʜ(v��h�T��Q>��C��(�Џ�*Δ��>
���^�)[G�^����|�F�`�=/��6q��P�:"����������;�7�`+�vC?��u���˳4�US��(} ��1�]0Gx֫F�`JB�S@��Ǔ_Ŝ��_�xs��P��561�6��S�6�C.��/�<e���a<)���J0����#�nΎ)+]��8U�-oZe�.򔿧 ��hrۮI��DA7%���r�Ҷ9���L�t�jؓ*�fWp�U3�����n^���s�O�͸���S?�
&���+o�Vo��Hj6|<;�U��8�?�9����Eb���;�8�y�,�Z�Xe<�����UP�ix��t�K��_� ���u5�by@�.vo^L @��.ח���l/+��ᖮ��=�Zfp"���5�.[���Ћ�t(�-&V��@�d��ү��?-�]
IC:);����QO>���b�S1'��)��?�Eљq���<��?� U��m^��-�r'`p$��t�����߬f4�6���Z:(�:��� $�E��{OUY"H���

[�?�����թO�^�0�w�2�ˈ�St�^�1c�I�>dZ��fi���Q�e,�0�S���fDYi;�[�!w�}��[Zz���û��̙�\��׮���ւr}�W% �����
�/���;B�����W�>���?�f�g�R�ݩ��<%���3�a�Q��r{x�e2�N�J�^�)m���	����X'�5@����ٖ.��7P�`9 xO�R��*V��i�v��v=��W�h��̀� (����@��B�����X%[su��x�0/��s�a�\*�f�u�*v-�h&��qi_���#}&��U��@H�T��0�k��y�{P.����(�r�������ђ�}�V<���6�E�|K��~�a�*U����$d�$�'4�O�Mn`(N#x�l�b
�I������?BU�p���ϒ�s�3�|H�@&s�,��{@��FL�i����)��]j����A��hp�뒝c;`���`W�C��K~�g��5��P���zڭ����PR5w�r�bՈ�2�������wx6v�0>��`f�!~H�&=���4\g�lu����wD"8d*p&���
O�.
�_�+f�#o9���O��4��I�R;AgvO��@�hŖ�-m�wm�$��Y֘k�v�� ��ERX�~�i��XWXd���q���<R������^�����<���-쨫�g/��cK�v���6����2�˥�w	O���\������H��Oݢ�r�l�C�OV����bJ��Q��Zn Gm9���a_����vc�̩Ժ�����r6�z�{�.E��o���4�`�L��v��T�՞��˫�^kiu	x�/4�:נ����!�Ɨ�SB����6n{��~t��[I���1brM�;z+�!����Ҩ�岀(e��c�~���ƫ���_7��3��n �o�"�9�!0@��aܵ�I�}B͞a�ɑ�y6S��$���>��n���.��PU�Cm5���
�M���t�������wtC�=��יD`W�i�Ĥ5@F���#���3�����©}@
�	k%`/Tn ^��[�?X�����FjRm� y�X�K��I�(X]������'�9�o�a�H��8��5�:V.|�Z�Q�Fxi�C��8#�����ׯ�EZ��àQ��Ɵ��ݹ��m.9�:�&*�!�=ڡ�Xe��#z��f��!F���p�Mw:H��3o�o{g~�u�4�:,�5�7����YR뛖�M�*��␥Փ����P���j�s�m_oW�HM�������4%c���1ivW�Y3r�@��/�\���1�2����FC��HO����0N%�ӧO����Y2�H�H�mJKlk/�K��3�˦�a�]_�d��� ��h�����B�ٷ�C܄�%��7h�y���N�Z^�GYe2�@�g�u�A����pL`�Ӗ��P(�̓t��	6i��c�hp���cݒ��Q��G�=�ZNmKg�T���������cR�u_aڼ����<A�~m�E� c=Y9Z|b��	ĵ�Bp7�zϖ��.�t_����!|���In+��]���E��(����&�m_����.~z��Pa@GU�Ɠ��ͻA:���}/�pIQ�$o�ȑ;`ݢ��ЋG^su-ZAAG�^���[���<�eqffF�'ǀ?]��$lƑ� ��yi_g/����g����ȣb�1��X���V��@���䚊�=؅Q
5��i�H��B3�_$��.����tBR��hE��O5�����\�@N��"'�&��*��+Ք�$�j���$��}��b�.���'�����?h�BY#���h`I.ddd�<¯�J�gU3�o_a��sCm]-����٩�^:)���kW�h�M�>O�#}�{ǒ$-���dݝI���}�p��I5n� #&*J���o�h�	lL���h��U�Z�#�-�l�ׄ�ߦ��H�_������9l�ї��֏�{d�M<av�^�aU@��`��V9���ҡ�)�I��7 G �֫�b�\*��2�}BZ-��= Jeʗ�?��2Ppvq�F#E�q����~��<�+05]�WD����nyD ����ɾ��'��ݵ0�T�R^<���Fn�ddb��c� �L��w�Y�6 �<G_bjF:���.�Ge�ϵ~��2��Pђp�|~�pkR���.��ڏ����QY�u�?o��K��&B�ӌT�7�T�H��ƿ��jh�e�n�-�+�ɞ�����Vj��y=�?Xb+W��Pيå����r��ӻ�bE��<�n����ԉ��ύ���S���B_����ѡ� 6%{����� 
j<�\X{�?g������֭�����Y�~�/
}kP����b�蠥�ŉ"�HJ5��K��0�������Α;�_vȌ�C}2@k.-t��'ۓp�.����F�~�H��������c�_I�t�GP������B`N���M����kK���\�,g�Di�0�$�<DE^C��Ji���3��Ju����DXe�mn��]á��=U��T�S.yy��������
Oߔ1�gh�U��.Ҙ��ƺT����`zqxIu	ؤ9M+��㬎�m�)	��~�v��~�s	��`xKO���
s].qj�����$�r�����ڠ�'
��B9���ԁ�ف�6V���ZJǉ�x:#��h����%�,��d�c�ܺ�ᠹ��&'8��(�+r��yM�D�4't�o*��#}���+��|�tg�5�}^��T?�������9$
�m�0�I�pi���	h��d���%]�R3�� :��K�V�h�*{ýK4W�z��U��wT�V>�<G�cd
b�O��Y�V���Չ=��S��Z�>	�Ĺvi?|��{��#�6s����B؋Ƶ���s�ק������;�%��͡N����?R���R�+�]�}��Յ/k,MZ��q���?x����`�2Tm�����i�h�W鎀Jر��]��!x	
��Ӳo���o�-͞a�TGO�h��_Y.��)zg�&��98XG���ɦ���#��z��h?��vj�hU��K���*����;ª,�;����{nŻ�|������s�����X�����Ns��=))I�ӌ(�$��jp{���o҄k
	򩏙��� H���}���c���+ڙP�ߔ
*���.�{�Rrzf�}��'����v��of�D�uG�0���uK��MLi���=�xE^� U��K�v��*}�O�E�l{{��B�<j#��[�87q��RNEC�RWQF�<zd2�֛p�@L��3nVci� Ήh�ģ�D_���u�JjPi3a����iX��\GBD�T�z�����ֲOVB�����͊�X�f2�F�x׍/�K&W�[��qP�����Q�]?O�\æ�w����㗍b�x�f�x8K�J}��=�Ayy��쫈�f��UsvECy�&�n�;Z�Vb��-�O�큁�W�y�>9Ն�D��D1&�QVH$rr��O�����	��<
�y�ڑD�5B��ȝ��ŶU�3ׯ_oޑ�ۼ�'�����1�Θ�3�����7;�V��I9h�M�����H�눛�_i_
tPX�IJ˽�ׅ���Y�g!��Ĉ&�����B�ypM��b�N� �̀QG������%���^@ N��xV�<�a��)��Qh,}�B:����'電�q��%��[/�+��
��j����62���+���=}��E��v���{�lcF��	��	�N�a�&LI�l�JJ:�Doo|��6�}�㔢��j7�34<&&Q�Kz��`��ξ��0ʝ{7 ������f����f
���vP`�]�f݋ �2�Y���٭*ϩs��wc*�; ?��=J���ȋ���r���\��5�#/Æ+3��A��9nZ|�*�X�P��'�RSd��=4�Z&��Q;rѭ�I���-�ˏeIC$oIjSR��=ڢ�, A��B��G����������G��^���s�p6����ڟk?'�2���b\1����R�9z_�Ҁ�����nA��G�R�ۗ@.�ܾt|X���n��k�POD�u�д��|DΗ�|���bl���xw�rK�@�1X������6�c��Z�ze���}��C�� 'ڍ�A[��^{�bk��j���F!�'e�r��"�!bPݺ�l7m��R����;��0v�,�]�`ft;8s�z�N8};^/���C�>V�X=)� TXT$��h2�GN�����P��'C��!�7ڗ�P�$
I�}~���=%�e�/��(�p��!�ü�!�w�gA�~P�ͯ"���SP�6�#,I�pK�,�b�G�dC�@H�|W���d�M��� g��i����C���t���,Ȭ��Y�
DT�B���_ZZJ��R�.�>[ ����9��l'?�r,�+��c��N�L;�7w�-�jQ�0��ˇ�yz�Kqx����t̨�Z~()$�w�F���Yt��X%:]&�/����}y<���~	ٳd��Rv���BIIB���	�L���D�Da0TvʚBƔ��)K~�=�������W��ɼ�Ϲ���뾎��o����^���o�����{�﫡��Q��vv�nȶ�0�܌����"���HHw#�y��u�=mg���wLW}6<����>���AP/습���q!u���2$�t��'_��,��>��3 ���źl�1���n������j�i��Q��+��p�t~X��re`����؍}�=���}}m���?~<��G��P\�����!�=����8����GN�|}��ɧ9>Y����@X ����qe�=��FT�W��ҋ�]$�m {�v�p0έ<5�XBda��4�&!��e�y��
�h����s��d���[腟�b�3{�l-�Px�f���'+9�:}����򔻻��v��"���N����R�Y7U�U\�ͤ��+�{�M���h�Tp�U2^�2c%�
�3�̬G�9�cr��$���m�qx<��>�[{�����3O��C9�vs{+�U[�?�y~��ѻ�%0O�i���{ U�YZ[����Ot矾t�xbb�5U�c��SG��8��faa��M*��?	v̾	���:�WI��t1 ��lz�2�4~����.���jj�����ݕp����$��tM�$ !]�\B�`k�5���~r�
82�Z�������+�y�n݂TT	ij^�!��?���J"�Tx�z����N��0�'&0�O~7U,#�X|M'i��h� S���� ��������ÜL��:)o��#J�j碢QU^=o<���&�v�ElO����m�A���*�|u�Aض�����S� @'��_���Rrjj<�q��*���d����Jq?���&��9z��M���2����S���볞��^]��^�8d�kdN"W<��,IA"��vf�pr��!1�Ìߵ �z��`��$���N��ey6e�N
A�c�}�9I�:�\�I\�)f���oH$[H\;<����w���Ť;w����`,��ۛ�C��n�����mK� �������X'�~�CT��(7(t�c@mDN���� 5-Xc�b��g���*��3�//z� ��3�C}ݏ~�sߖ1��	����/UF�����S�&K�Ig��v���}�@J�,��2^ HN࿣������O$?����X�`/&�Fu���>tjC�Py�#��顁Ǿ��7r��]�m�4��J�*�l�H�]X�����{�x{�B~�lB:��+�F�-�NH����%1I�hVB��)ڄ��}�Ԍ���@�n���U��|��%�N�y���4�'���/����(155�W��{؉�Y�V|��j���A���՘��K涑��x7O&z��K#��[qi��_��EK�rF	�lBz�5	���w+��*X���BS���?�-(��Z0_�3gK3 �X�O�<ۅ�X��^��J�dU��h�!˳�B����9b��7'��sϯ�D{(z-������u7��v�-�Jy1�t�&ͤU��1�rR�߈�TCZ�)�	-_l̵�5{Nz	V���+����q/�S��ts4���ˏ��2=Mo�;��ж^�������pY�ç�f_Q��t6���[�9r�_���Dʝ��!�$$�>�ۗ���m����SN<V�c��s�y��?U���Z��n�F��+Gvt<�p�1��tBjH�v'` �i*If2���xO;�e�nC��p��G
a�Y[�^��r�a�����$���./N�_��ԯ�I�>�=b�t�C���έ�Vh|&�W��*�s�2�t�;��u��{L�&��E� 0�Y�EK/�޻�qL�a՟�e��&��4H-<�D����[~���6�m���q�e��!_14�[xֶ�ȭ���.,�@�����nXw�>��A�w�]��I�R����~������q��U���۾l|����G��z���m��X�-�BZ��>?sT�о�Ƥ���t1{��X�K$�=H%¼{=�F�0>���m�,v4��B2 �R[O���ھ9H2�o<)!���]���o?�ӧ�N�-�<AvN�/�-��PP���q�����_�M�`Y�u=ȭkU7��`(u�=/��	H*�{kf��2K��T��ImfT��LS~K݌1gO�I��nS�j=AZx�sP֦\���B:��&q�0�^�����Q�4�О>����Ks���w�1�͑Tp
�[>ײ���H��{_��~_'��>85�^/��!�ʥ)�Ї��L��dٲ����%ev�6Ny�Dו���������ę�r��:��[���$BI��~�Cg�ƚ�<y�y9���W;{������{W,��b�ZC�Vn{M�;T�������B�(Q�����pQ�#y�ؐ�=q���~��D�*:���*�7��S��Ѱ�W��� �ⵃ(���0��s�Θ`qB5 u�ک�K֎��/���ǽzu��L��hWb�{W����s]CC�hD{�&Q5���B�~�(��`�2�l���~�j�0{w�ހ�bF���iEhfV�a�<����g�A9=�,�KY�J1�,���������݌ ������+���kw��{�e�_���/"#u�8�{�~4�O'���g�j�$��m���I !����q]1��Qt�iv��x����������i�~{t�����a��\��� �[�����<��~�h�����ҿz�\��r���^J���Ծ��v։�P����V���{���G���mY�TȼӤK�鲡*h�wQ?�H�Ks|�<�֐B��Ue��t�7[�Z�/H�(loA/�4�-+�����]=}�x�>|lvC���sݽ��� :���K�i't��ގۯ�Q��� {��U�1֐�dGQ)R�=D��o���WޣzŮ��_�C�(�R8��*iӺ����I���s|�c�N��t`t��.������T����O��L �G��GS�� j�^�T2�S�Hmie��<��x�B���
n���(���@zy�M �{j�k�W"�u��H�z�݃=�1�h� ���Aź0�Q�$��Ր����W�k㑵�R�gϞտ���`<��Ȓ�&!��5
,���m��HN:򪲸L%����K)H�=���H��'�/H=�C�O��%��	1��s��j��_�ۈ�r�� 4��;և7�Gq���������A3����� �|Dm�o�6碑 ���A��9�$�o�s����c��QPC$p�)F"c�}C�nͱ����R�1q���㌼>\9���%]U!&H0}E^B�g�_�/�����Z"���L���t0 �E���kwxq����O-²��HC^*)/����p�Vh2d�#�9��||ԝ�������Z<� ���9�>���=٤W�.��0��a	�OX��^�λ�$�,��@z�)��Ra�-���}�k�j�3e����i��S�y,ͻB��#gu\G��� �A-
Ya�DVZ���Cs$c��F��j�w�!��F6a5-4����"�Y4��J�ɂb!���y��Y�7W΢��py���r	�|#�b���.�I�fX궓ȣCQ���#��I��}��͛���?:���Ê
�e?!��Ȝ}��~r4�1j@����^z�Z�����
N����*���à�hv���:�V�Ε�Y�AJq����xj~�����p�
�kq����ha��a�pss�|�����ccy �.>D�L�ߋ!�<�,T:�I�x
���Z��d��zV�A:͙�֪�`���ߢ�xVNDon������������3��Uw�|,~=���p��.e�Z��O�M���ϗAg<��NMO{����ݱ�������vBBɩ�yhh��-B�������,)�p��=_/s���Bȯ�ʘ��<[�.3�x69� �E�6��]�M�e:s����QaϞ� �=,*�L��W
��1OZ巼��-�@8�ߔBw,�?���PR"�[橁
JΧ-	P���{jH z=8>�:{QA�z2�������q���R�ޖ��C��v:]��<�r��
�5���%��>�A	���=�ԮS)�v�[g|_j���}��4��!�x�G{��oߪZ;:�wGdt�D �BU��'������CS�gV��p�d	�Ւ�4��N�+ij��B����� ����o���^�1P#ջ:Ó`;�!주}�2���z�s_�X��	0G�?�
����R�HQ��n
A;m�gZ|F�c�RU�L<g�/I&S%��.�{U���ٿ�Z�v�2���l�l����#x@�C��v.���@����_\~=Ԝ7�K�M3g����hm��,����3���Z��v��X�o_"��X=��J���c��x���Q��-�+�tغ٥/'Ծ���������w(�h

���
���z��g�		i�9�$ymo�Qn2<B���'c�������^����%S��r�-o���;]U�^tg���6S$���
����sW�:�_�a�c�{!��~�
�I��e_}'�x\����ݭO���u=}�g`k�cxȿ$����= �ɢ�Z2��<���`՗��C�YC�tF3X�m��9^=n
b��5yT���^�LE�\=#-濫qx�yw���hqe��V�;#�Κq�dp>�rǔQ��:J�av�ޚx��i@����>҉wVE1�-�|�5/W��}���D����4��/3�Z�y��b�,�jfs2_��a��<�6ȧNM���b$��ʩO��D�q
TWe�<YxQ^�ԯeU��g�Òrł��_�QX��U�����/Z��b;���8�
��\�����$�H�*&��ӈ��m/C�<�'QY��Lc��2%���"�!�>��x���f`.c�"ِK�My�i
�`��eb��74�a���!^X������*'p�6a4�`n��L�Sg����|L�s���G3�(+�T��.#n��!g��W�v�C��z�ƹ�q��s�r��%�,��Ac�^Q�pf
��e���΂4`����kM��ϗ����뱩v������n��&}o�薴��g��9��{v����ܲm�jؿ��M���]�s8���k���wH�Q�c]��	�2�e��-�`\�����
��I��ޣ�����I��3Q����~��zPPU��0#d���I��u����v���Nb�bZK";�r��A0��w
Z�[�<��q���~_G��ሺ���G*�A�_�F����=`����d~-t�~�|�KY e/',O�'�H(�@��3W�g�/���R�b�� ��%� ��lvHoU��urhM\0�X�C������� &Fm��oW@8�řd��Kݺ����D�:-��K��qVUZ�w�i���D���+�m\hx5헲U�j��/u+�fpG��puAL�d�-/Kh�m�+��AKඦɗg�j(��h9�@DS0ߒL �T�-w$��+���K�U�쯾̳���p����G��?썊�U�L�e|��7BE(�E,��N��̖��
����P-���%89@�\��!�M�72M����EdAÒI*�<ʟò$Y.�_d^~?Sۄ�.9C�͗T��`3�����b�ǂ�ͬ�w��^P�F��� �@��4�G
}l��o��O�p�Q�[���H�W��C�ϑ�r=���}�z�{�%]V4M����n��T?�����fݾ�g��Q�_:�� B{���C�ߎ��]��Yb������l��%-Z�UT>HI�5��nh�$�͝cy���X�����7+��u]�*&8�+�V�1%z�ZUʧ�p�	��I3Y�)���3S�q�*��M%踸��sP2X?'x��s�;3\�o�[�	c�K�$h��oS0���S(��]�=�%�t��:�����9�E�`AC�x�r��@��@Ё����lv]�sr�Qu����z����>f��T���'!�t�N�#-�G�璭����	8.ݡ��,��D����ǝE�D�<M6���N(W6�G�Ü7胄�$vA�a�XqN4�8��ݶ��n��;����r$k�)f���4x�-��Ϛ��zD�U~9�������;;�Q�!{���:A��m��.7�MzRM6`��2����Gr��ڋ�k��6��Ɯ�͟� c���#%E��*# ��+YT�L�'���bIP����_���:�_�+j}����2�������Mݝ ���ܞ�A��;�U��i���j���=;�J>���e�������Ȑ쥷���޸z�����0^n��A�_ţ��`�j�l*��RpZ�$�/���[�u�h
���#ǇuR�Y�_�C�8
U@9�ߵ�|�VG��:rd�6˯
�������x��#W

���z���^i����ƣ(���4f[6�/|��P���c��L�u�@������cx4^��D$)�lHs����gW_^����k���[n�w�����������ia5�
	�wA!�r�a��3e��yck��U}�+U��FI���_�b����%��P��a�Xu-K��(�7/�������:!�0���R�����覎Q����ڿt���57}�6��:�=����s��n��*ݪ�+���,�zK���M�x��Ao�xG&�M� �+3���=]���Fk������Oo��4�������� �lh�`Bz4[��١� ��A���1��4� w�m�%<[��_)<��^{K���>��f�t��n��,	ule��\��&#m��9�n��VXW�x�A�����yRM:Ww;r�d��	ߚM�h8nH5���#�8����Q��Y+��TEiO���o��+c=����BT�oF�Sr��{B����	�w��c���1�u�&mz����i"0QN�dΒ�z�M�vYJ2u�NA[
�s��������������H�9�t���H/��m�L�3D�M5�qH]�GDvR��BJN��Nd���yc��a>�"�V�) C��eo���LO~�V�y_�A�g�N�֐T+d��i��0�ϼʝ��5fؖ�,5p�R�i���w��}|�5\����v��hfVd�bJQ����}:d��$u<I4z�����_A�k�T	w=���7��H\����*�	�þ�(��o�.H������C��Jq@��҄�@:R�7��dɗ1
W��%�+�x�	�g���6������]��\C۶�D����|��g`���4=uu+ǇO_d2��P�T�z�g�l�e��2Ś�zʡ��e�$P�9*�x9 =_����9�Vۉl#� ��o���{h�2uh'�kk�.%\Ɋv�$�r?��� �#t�?�6���M���h���0��M�s�#�� �Y:�Y�-3ņ��A� ��HoT�2-�RPB�9��,����51����.J&o' G��f���l������9�v-Ȳ��&�D�X�s"�{����(��V����m3=P����U����?����.9#|G\'���o�􍬭bu(!�!f��ut�CI�|y6����l���X#Z�K�x�&x�H�w����{y��JI��t���������p��ȕE�/C�H�����5�Ȃ��:��nS�m��� ��H�e���U�Y��^�Q^�ci�&d5�A��3ଘ?����_]����N����)]"w�˖�֤ d��|׉D��bdL��F�ʊ_��d���nȿ�qЊ�F�x�Id{w���|�����60�Z�`�'a�̛���M$lQ��5T[*b���a��  �f֡0�AD���{i���׬��ET�+;��
i �#���M�f��= ���z�/۩��'Swѕ1{Xi�bD���L�c~M1}g�J�<L�9 +6Q�*�Ƈ��4�>��\$��s5K��
`�ZbT�/1	�%[Ξ4���ࠥT,�"4��.�s�[����H$�Q���v���H���J�8�|���v��Mt���xbT˺ ��?�~�:hq(�����&h�:A4v�&��s6C�`9B���-���!��;�a���n!�b�a�h0�q�.�_uz���}��V�)�Y�t  6�F�s}s���6���[�����P	,s�
ҫ�@�<yS�΅0�U�u��� 
��֗��'����>��1!%�N[gA�h���uS(D 4��gy8=��9Q�O�/�o���V��gN���Rue�Nz����U]u�8��H�&J(�@�Y���]ηÎ�����܇: '|YLzq�������g�NynY��m�#��s���i��i�7���C�n��Է�d~XGD��A�0P��sV��[(�^�h�9�V�
��-ϟ���:���D^~��JC�>���r��:�a���F����i�Q)BY�S6o���Z���Iha�㮋�3�~��+�~{���GA����Z����JƉoW�O�8�vn�W�~���������}8������ �x��q#(]��̩�z��x}�`h��h��RG ������f���ȗ	���­��}z}���w�$NMO?_Yy�����)
�Y{;�؏'mC(���$R��o|�[>|��w��'j��p�z+��2/?s�����$Y+��{��6�$=��-�Y�����`M�lt ������#��Ne�I�;�IDSNC�
r�,++cY�.-�S��M�@=̊K�����G� k$�a����mg3��5�N"%�]B��$A����1kRd�VlXPI����������6 �aq2v�.�nq�4��g]H�׵�@GY��t:s�ԙ3Ff�js��������7�-��2񥥥�����2�W�����o��/� ��褜"X7_4%y��1���$ b�f*�i�@MVT��ތ�/��}���kuhmk3�43��xDEE�@ş�qI�@ P�ɬ�[�L6�Q����~g �4u2&�`��� �fi\��a^�é~�p� �l�2s�+Y$
�`�|�EF� �K��24vv$3����K�j��E��>8�|�)f��#�H���cUV'N�?x��_��H�Q���udP����X��9*��t�̮I��oK�p����o�4b߲�V�N�-#�*{���9 ���1ӯ��_��~�c�����+O��{u��㏥RR�L�3��%m{ie5��O@M�g ��%���̲��9�,��	lf�aXi	�&�����֠�?l�9:@�P1�{�(7�d\QY����H@��pM��.�]}u5�d�+W�)���q��.Q(�bR�%�fc��<A��+���Z�s1x�&�Y��P�>�����F����w�_eȏ��~$�lM���.����A3�t��i===#oWW���[t˝�M���ԋԺ�s�i񉍏��X�m=�~�6�rN���Vgk�u�W���Ӛ��c�OV�����u`׌�9"�����D\g���B��S� lv������V
_������9e����)�&eSq?�IQ�MD���D�����$)��䲪%
�SB��8:y�>*3wK��L�2XÇ�<�	@Eϙx3�Z����!�Q���5@������u� ���fꐴ���)��ߣ���ƴ�����P����$�s�V�,��p����C����3��R�
ֵ����� ��ğ.%���� ���*���T?����x�s�B��8B&�+�.s޷<Զ�������,1��=�b�K�n�L����5�W4�w�q]ָ%��xP�A{�����#mg�H}?����9
�x���>6���3�v�i�e<\����3��7�����"������\��Z��ݽ������c;�|�CKsb {���X�H>�<���@u>�:��ou�L�2&U����W,c%�fgK 3C���OV�.Q�q����[��Q���
TgO�T�5(�n��'�A&qa0�w@sq߭ћhȎ����D����F��㒓��/A�����I���\O�GԈ����P��}����ي.7����-����΢�( �?�w~Qh�U9s���(�/�#\U��&vWq�^��'�+����вVW�..��dS졘��#bh�~��ig�hF���{8PMbOqg���c ,s$�iΐ�vsݗCֻ�R8K�:^'UB.	���ݍ�ޡz�r���A��c�6[b������㵌��oV����t�����G�3���t����:�]��JYd��C��v��I�������?�*��j
\�g����e��o�K�~MP�G�چ �0��[dr9�?#X�X1�:C�ߥ[h\���O.G�8�fZ�2��+�I������+9܏�R(�qը�?[����P��1)�(�������D*�v��x,�}�1-�D�<����&�<V�����]��F�ǁY2�?�$Z)�Id�~p�7o&��VV�$Toaf⽆.ݵF��t/��|���9@�_y/�/�T|��-uoP�c�U��Ox~�(��u0Et�(!����qy���V�ǻ@;� ��r���B���e<s�����=�����ߍ��"S���+z8��YWWS�jo��qg�Cfq��=��*��I+���D���ڸmn��W�B�U>�PX�ß�U1��z�u���bw�
���'�>=�_���KY5q�%V�����nw�t��|`xi\rd��.��딬�E�J&��{��!�C��;22�t8-�r^������ҷ��r�Z}��i�;����U��I�VC>�h" ��π.�N6P����U�21��~�a��G8�:_��we�vh�T����������5y�� ��.���H3 :�[6Td�7fCІ�?��q�0�6�m�l��@���I�� �+��HuԞ��|�H"	�sm�v1s ��h.��{M��h<ׂt�7��e��V��Gs�����<u��y�P���~���<�f��f��棬�����?W�����r��
�i�~x�ӄ�}�%s9�)P�3��s����J>䲚���� KA�2!��L�/2@A9����dpO�:-��D	���n�Qg[C/̛vi?'e젺d�n��$��v�޽�����`{��c�7{;�F7�6�м�#)��b�R9�֪��*�J��6nLё��)_�p��}b�WFN8�RF�b�Q�)��wN�ps��`,G���ݿxA��D����o�*��(�@B��4��j4��C�����]ħ� M����*9��|KW� *Yp�����*�<a����׳rv@�G����o_�,[��<�o���W�Ve�껋X�>"�=Bћ��8����fL�+�"<YmU}�}�s�7���̬�9�� p	ŕ�Wń�f�d1^C����*k�OJ�W���,�`�D���q�׺�sY%YɗA��������d�v�n�EJ4]���3��0c��nOU&��4Y݌�x�`��&)'i��� ���o�E�'^�r@�4�]~����۹.���H�怗�缪���-D1h���a�X�3k�H������#�#N��+秧�ə��h�����Ѱq�`{yC��$����-��GP�A��������]�Ň��9����ɘ"�'~[_LYz��+�5��ēk��Z�*�8�?��g�����J�����w���'q?�����z�x�+�B�XE�v�W�4yB�.�u0��v���7��:��)��Ճ��H���>-o�ʈ�=�7b��σ�OX�չ�`]Ƹ�Vj��;��M��J�D;I,r��v�k��|k�7�3��r諗��-��toՓ��]�O��p�r���7o2��%@">��[����)ïH�w:����벟�h�e�G�͑T<�9P�����ڱ4N���i4	
4 :�j���(�l�X�Vξ�6�
��a�ֳ"+k�M2Y�|��I�hnM�����z�M.�;=��A%F?��CeܦL�$�1�Tm���n����:y	>w@ ��b�{ϖ�u��7y�<�!;\�V��g)(��mj�NQ�3+����쩰Ql�������3N~���&������Ո�;��*`�AP!l#�Pm��,�_�:�ʆ.[nF�8��J|��_���/�<�Ռ��������lکb�q�	^y�H���9˺�wL��(��^fa����ZI�x�5�$���������M	�;
�O�}�]��U����g�e99��o��z�r�<�˽�ڋ&�_�ԋ�S�GJ���Ƕ����x�G��ۙ�8S�2 r"������?dqY�_5��L�(*/�?_~���wU6�`���,j�H��[�k� YTT]]=v9�?�a�8L��8�D�����6��c�:���cZ�4��*ͣ��D�PT�ﲝ�4�Q`�Z�䮛��i��2eM�����%�ND��b46�F"�â������G�{�9����X�<�=�}�R��H9܅)2tg�jJ�J���(�����E���3-L
 �>Mp�e�&�b��Ϋ�~����E���v_W��?���U�9d���Xc��m��Jp&�W��"���"�h�Y�=�&e<����5�h�w7��G�i�����eo�_
�J\O=`e�9��O��c3�-�H���������IAm�{�.�t3��������GjH�� 
��k:���b�,��C����#�y	�����o!���4}Kܣ���Z[��F!�cc�����O�,ң6��r�2�B�KM��6��6��ڰ��	v~������xs������#����,�	p�Z���4��/q��y�����e����t�wW�~�迊 ���n�ǂS���ڕ��C��8�$��$oq<���z��.���J+���`����� H$��gH5FKJ���Z�*�Y���4,3��'�m$���6%3Ju�k�
��.�'eff~Q�j8Գ��.��_.dyO�r�����m��*�[.$5@��!$�^e
��$�u6�E�1���B9��9|@>�$����@)���[��aU�լ�$8凅��khh��z�s�!r�M���ʹ'�@2��_z�S�PIe���f%���ʒ�>�[܂X�ϳGEɽ�!�3k~�p�h?����.�z�w�������:B�IG�ы�TW"z8���]^�W;��sY��{]K I��ysEh8v��Hq��e�ǘ���w^1D��C�.��̜���ۄ�4���H��ڝx�vڈ��;�`���"$ES(րѲ�Z*��<���Ӥ!@��5q�59WA�k�L>D�˝q�!6�K��|,�"���o�ʬ0|Z��G�������;K�]�B�!�5��p���qGunr����΀*'���x��ʤ��������o�;<��T�w$�7'+9�7~�*��?K' ; �x䔍��bO�{�M��qA���Cn����t/}r��Ӈ� >`�hch��	?>�B�䬿K�%��&�]��,4���hΫs-w,�On>�[ʽ;�׃�i��ֳ!�l3�&h����͈H�K;�9p˿JUf� <�	�@�bN)�Vŧp-V�
���Ը(�ў�]i�>�)�<Q��~ڐ�P����Ve�k2..��]����s^=`F[p�lK�Orw�� B�m�#Rp�Оh*�h�"�#�zx./h4qY���'2,��gj}�R��b?�j��,kI��o
��i�8��L*D�Յ�#��q��#���ʎU��X9#�[�����0 	�-�s���W�Q��G���fn ��v쀢�d��h�/-����-'�!��$4V]E��?`t
��S�<�����j����Ӝvw�B��/���!�� ��k@�(a:�w�v���F֩�n�B�|yM��4��n7G+���[��?o�n����M�u�����ՈD���j���T莹v������Ï�~}�^qK�j,�ːNYZ�z���5�z�rɈ��@�-W�e�(��t
�M�����x��
]G"�@6��垜�D!�D&'��O=	�K���:�i
Ũc_� Ͷͣ���Z�Hp���[�WX)�l�>(�Y6��PC�Ъۗ������	Zv:�Ñ�ީ9o���Ù���$��7��s����%XlN����F�$�#�$�1H�����Q�d,$ԁ��z�����[Rba��"�RMs/_&T-���
�Ҋ��;�G�#)E�rcՙD���M	��YLck�`+˟zTN�+��܅�G<Ln�!�V����B��)rvU�LLL���A�^T����5��Αv C�v
��q�ƍ%�)��^�T�XR��6�F�h��o�Gr����PE�h��U�LF�����؝������T�����>85-9HMӉ����%�F��_��^�nQ�Z�i�3r�Mn�L ����U��qʼ�;[O�Ͱ�+Sӫ�c����.����U�Cb�u��i]��:،/�Y�z�bȕ�h�b�1�fT�5� ���|��~P02��y�Ϫ׻[
*��J��P����P�T�����J,yyC�zc����l�ҎŎ?m]5�]�E�k��N"�Ծm3{}٭���tuE%�ύ�+Ch�Sj�8�*H���g�h{t}#��y���kc��,h��t!�	�޸�1f=��"M���~a�[nl8���I��Hq-�hxG�g��N�M��V�u_��>���B�_����W��U-��i����e������������w�E���F�jv�{88d3�8/��3��[sc���h���8}B�J����c���$D��)����"u���Q#3,E_k��z:��VǴ��"���~%�яq�yܭ9�|U�!���Q�n�S�.}�����~PoB9֟�D�T4BUδ�?ꉙeE�r�	�\"M����7����-֎#�ߒ+���C�z�&@,9'��"�;���7?g����� L���qlZ���W�ˎ�+/l\�����%�̥�T��/��R���6�|a�H���8�����R���ƈ;[��i"M��/[g<<�g�ӈ�	.0�*�E�-�7r��Q/V�0Ư�A���f#�?e���#��Ɛ\ʂ�ax�Ϡ��w���Zq����vg�"�� 	W�uf|8��]E�ܣ`Y8���-��	�ƍzX�+��@��é$$*�
��Z�T���j�+w%�^3wM�F h��؈���w�HAo�ë���_b�p����kPb^V���]�p&[8�OpH}Gh�{F�p A}PN���bL��?)�̥g�� q��x�ׯ����Wq���>�Z����t,dX���疢=T�51L�ӥz� ��H��!Gc	m�)Vg���B�;g���'�� ֨�6�b}v�W�7��k$J�.���� �e6�X�o�����B�s��^�Of�}L͍����I}��W�(a_����������:� "&��]�<�y_�F볓�c��
.��-0K���Lw7�!I&2	�_��2}��4�^t��6�%�"�|9��m!To�1���~ FH;���!�of�ڻU�EZ��zqڭ�U ������/Je%��Ifly�Z���@�9v:lS����SIҍm]rz���b���
ѰK��e¯�wd�\0�<�*p�]Ver��)II7�X�^𜼬_�����q����&��ǈI[ h�e#+��(�C���*A�.�@��m/C��w�t=Jaҩ��;�%im'�������ҧ�751���I����e%��qݪUO���H{Æ������]��
���^��^�̤��ra/aW+�GK�o6>&\���)��VtL��7/n�A]�J��Btq�F���b�G��ѣ��*����H��?C���䣺vN%SV���aI�'�M�V�A�S�����6v�	T�[,���3�Ӥ��BCmm����"X��/~)�O�P�� �%����qh!w
���W?ɭ�a�߄�gȼ%����ޜ�Ͻ�
s�?��."E���E�?��5\<�|��.�x	'ç���+��QK�~F���c�wR�3�:T�6 5�\KT�����>�w����%�4\*�=�yzmp��c��l9�" ���~�$A�˗"��Т�����"{z<|���jX��FD�Ne�`��C@Pa��'|����_�_�[��r�����㫺7���y_,�:sh�>ɲ��T�d�\<�|s��+"ЇM�鹸rW��H���Pݨp��&�[�]{�P�_@�
w.L������Wfb�;����=>@Ɛ�fow����<v���N�f�.±Ǐ_i*�h�3�އ�?�?Č�aU\�#O[�D}
�[~�qO���-����>A�RSk{���8����
`g�jiْ��Q��q�����0���o;�Z[Şoy��{�VP}'v����[=	�;�73�1�E���tU���Uu*��VyT����=_D�d� ޜ���}D4�b�M�(�9۟�d3�u��Օ��'~�Ӈ)�g/7n��OKO��z��މ
���Y�XY�"S(/(����������$v�d9ze���u�ͬ�_�l��[+�{��$�s����0�[�x�d�G��j|q����+��S�2M:�JGMPUe����lpǹ������B~�s"�� ]Vͪ?x޼�����.;V�A�p�bo@�D&�K��M����V48xee��j��������Z���ϒ|fM�C*��Y:(j� ���$��Q#��\D�R�NǞ��"����A\?ہ�]OE��j�vT�ȸ\UD��,9�D�%��b���W�n��R�^��<(���>M��&��Fǫ���_^Z��q�����ꊜ�߷$@�;��-��l%9��)�7�rw��s�g`���[�~5 Y��龎ɩ:b%bTUz��q}#N�����E7��|58-%�Ϯ��\�w��]R�{ulve��Ü��酉�cG�d������� �44r1��ѽ�/^En��#]G�	֡.��=�K̽��S;BD2�0�l!�����,Cy:������k}4rMUr�sH��c�_`GkP�VDԛ�}P
�ԕ������|�H���>F����s�'�W��ũL�_�y�5{�U1'�GSz�E��.Nv�$�)�W���ك�
q�.n�`�1�6�b��}�� �}^�%�;~�^g}6ɏ�X�M;����i�*��97?YY�ۋ�o/s�s:�3}h�����W��}T�=S�{}�,W��E\-��A�]�ݪ'���[�q��@�$�BW���6��杦r��ݺW��29��x�'O�������b����#���qMP�o`˹����zZ�B�Ȭ�����+Ƈ���Wح)L���.��K*<��u��#�]K"o���pP@X6�cLjgͶ����J�
�MH2����XM7Ț��y|��WtYy�3Wv��ɒ��7��|�Ff�_���������>� -�������o�!.��]_�.��B�u=��Zn��|�=H$3�2!}cIv�^�S߻�J��J+�m����9m�����t������_��ж*�`��|�΁���|\�;�᪎hXL�U���CE�$�FܼF�z	FJ�vn�W��Ĥ�f�m��~3��W9�4l�%��\�9��d��(��'�F�<��{;�cږǵW�O���֑�
Cy�T��j��;���c�XB�	��[ԍ�����P�������,��Ou��֢�E<���^B9se1�aay�$fI5P���2�j�F��E�jhjނ,�Kۣ��-�Ѯr�%�ONs�v�tj>a���t��y�8̢�v��[s�0͠F����5
!z���TX��;�����j	R�U9������M��.C�����O��h-M)�i�-�^h���G(���,�s%4?G�|�RWd�@�<����/3����������� g�ED�Yξɢv'G�����s'�>8��#+�+Oa�U�FPxVE8|����U����[���,ϓOx/Ξ�:�K�}��o�w��=�����.W"��� R��sV�&�F��f�z*�P�����Oڋ P�����0� ��x�,
ϳ?$i5�*86�ῢDL������]�q���E�I�e�0���.���S��x�&s�>w;\�,�8#�/�RX�!8�O�D_>�ϒ�9�\��(��K�A}�"�#�u��������uqrS��D�Yn�+l�g���p뾉���7<	Qpn@��H/�b�ni�BX4�`��F8��:n��A!�(f;du�v����ijPJ�/���������/�uo޼��9}(���7&�h����}��<W���^&�w�UN#t���n2X��Ŏx|M-s����&Xװ���775ҌKn�X�y5���h5F_�z�C())9"eI*�<�Z��D�?�-)������k7���@_ی"T�0���(w��%�8o�{,{0C�YSo���4���9���ҿ���t�X�z���}�A����8Cƿ}���{�@���}�H�Q��5{ei���i�dْɒ!"��F�}+I��24��ʾ3F�B���~�=�>�?�����<��u��\�9�9�&:�r���#Ko��Ƥ��Ȝ�b����_�#J������/�j��z߀��M��-��\H��Sn�ô�X����v�������źe�*
�B{�j\�i����Ds�d�*��ў!����d�p�6I&�!���WMk�Ʌ.+�@Gvs��0�ñ�j̃G���Ȩ4��-,ؽ>�1o����)��X&�k!q$���'�_�?~�{{��ˉ�h�,A �}�W���U�J�)k���>��E.��6u]B%��C�w�E��B
���e��Q����8��~�PM���9�⟞B�m���R)ھMˡ���������k2F�X���{��P*���� � �ƺ��:�6rÄ�ePѽJc���㠦:x.��OZ�L�A�a�X�^��xT���*�?�`a_�A�R��&MXS���\(�l���ƫާ�\���u7��2�8F{�wiԈ�<��ca�A���X�S
̃ԋ�>��)��~�.�g��~����1��j�K��
��g_�Cz�� �����5�������Ô6f�T3���,�0�����.��k��,Ptgm��m,��.8?��%"԰n��'����sl�1>!���C�K��-��1��茂>�����S��X��9���}�j��f�Jq�1��s��������&A#���`�b��Y�d�M.��˝Ty	]1Pi�_,EY�m����{�����V��Ű"\���e�|z�����#B�#�?E��~rd�ی���2��9�%0�j����=��ϵ�qb�ApCT���̭ ���{r���lW�\��L�� 3h�j}0���˓�"&���UGĒ�6�8:�o��`���Ns����I2M�rn]���|Z���<wGX����$��!n)��P��J�UfR��kàǾ�4��Q�S�ڿ}���+�a�y;z��w	����%���x{_���VR�"ΐ�@��4����,f�����/���7�RVy�E���G�W�J0�;�<�z����C�`7�֟�	��H�Ȥ$��j��k��aL{�+f�^K+e�v<�GIZq�~Tx��qǎ��Uv�'�*c�q�F�u�޸�Ƒ}��ދD^�H��E��V��8�ܐ�fc�@�탲���P����� t�|IF\Z�f��M��Eze�(%��+��9i�稹�ȱ{��! �c�];ݐ[3����RYS�+wNy3���BH��4���[�ؘ�Fc���<{oT�daa�7L;>L���rݶ(M���=k��C;�-��a���|��,�&�<�5�l����u����=���aV�څ_��m�����B�e��a]O����~��)N8�յ����1��AT�G���h�=v����
_������ܟ ��bS�ʬPq��+l�u}��y�E�7�RF$g�MH��Ū@2�l)u<C6C�@ݺZjR�� � �"hq�D,N|H�]<��,�DG����]�FʨlN����=b����+���K'�')��>��<=t�Y��n�m?� ��l"��xbYپ�H���P��W����}�	A��G�h��� ܒ\���ϞϬ����~S���JV�q�!��u.���d�+:�s�l�aW��.�B�-����6� ����^�x��|��辩���v��"�����Qm��w�ZXؔ�q��l�'B�	�Q쑓�����#
mQ��-�;W���+��kM3.��xD7&X̑���x?"U\�>�$��� ec���#���)i"t������O�6`e����y�[�Î�#pdG�Jq�>SrHnA���2�z=@���D�)12��V���G�Y&�[�������i�dl��2=���N�ܯ�˓��@:�n�@+�L~`�@�PW��H���H��TzRA�I=��a'U������d%�D&�_3.	��v�*� m��CJ�؉���J��m�'��>�b	R��ذ �"��\�;�ݶK7�]���}�'������bEb�vI�7�ז��R�b�\����׍;�G'U�f�������38;���ٿe�(4i!�(;��y�ڽ7�|R����X.�a��ƭ�f�gM1���ꊙ)z���5����ގRC?��J��L�Z�*w�C3&�Xŀ�v��B����"�lFo	Z(s��_* &&���
�j|�D���qg�{B�u��V̆�-��лM %�[��f�ap�2v��I��tv�>�;e�%�n�f����i�PK��4�N����=���Rqx��F��[�HܓX.[a3�r����:v[�ߒQ�FD�?��@v���*�R�XF�o��b��V�...�=9���ھܡ:�v�[	ӻ_ަ���@�9)plOjªn[K�q�27������BVhn7{��`����ӭ_����O5��*��2����u��H%O�9���8�dt�hI�Y<t��3¶H|���1X�H�H|�ײr7V'u�<؅)���ʛi=P�̲C��LbE����"&�A$�G�-��:;��Jm�6p���4�` �|�I5�]���'Ԝ��Er�!�����6�l� xO݆�K����[����u�}BtTZڽ���)6?_��>.��_F_ۿ���P�<0��Q;q�)"�eɴ1|r��X����F����0�W�{�4(E� ����5�ޏ��w����w���`�.�$ھ��7;���T��F���vMA%d�J+x�U?��@J�~�����N�|��E�z�t5�'W0�8�;|���M)��-_�]��>���_w0�����	���miiQ��dk������5�9%p�ҏbIH]�{�i-F�Sq_��BV�> �mVʖۄY�J�]��J�^~�׺��t��`	��@xs��;���.9�~�x�ck�{w(��Q���{�k���LNX�EwZ����k|����c�#R�r�O��?��C"�^���0�	%sG����QOXx�(�N.\�gȋF�m#TH��W�KLN� 8O�|�h�ӳ�N��=�_����zL�!�0{)�f&3Q�2��*Tb�������i���T���H���f��K<�`>())y���th�?�׵˒H��'Ĩe���͓4�[qƌ��~�¾ty�,R ����,�Y`p!�V�}�%�ס6��ԛn�Zh.�d�,^�;g�%������}�ꆥ�}��*���{t��j�8��$ �(�ó�b��U������>��VB+�9W�IX3��Ej�p�h٥�O{c�� 5��/�4��squ.-I���[8u����~���+'���&�S͚�l>���t�0�����vk�V�&%� ]����֌���X�(^].t_d�F��=�Ь�х�X����%s	��?�￈뻝z����	�c΄$Bg}���AA�A���8��1�t�%)3*���y�8�����Ѡ}����w})[4���`�	�0,���
���gBwv�a�vjikO �a!���bjh�t�*��8��u�u��s��z߅m@}�cB<�=Q�	�<��Ĺ���!�;@�T��$r� ������D������펟�wL�#T��īM������U���KiD�C�2}'�"��r�R�Rf_�gN�	������Q�»@��e�����H�m��ssgyN�y�65�ᒣIɴ�aB�:]t�8n<fF7����H�C�-o����D���!U�-&��8[�xR�@��{�h�v�->E�����sf搾܈�Y����@� � ��0�nR �%~I�2����s��h��9~�B�J��e��t�OH��D~{���!�c�C�޽ѫK�@NNNѳgZJ�M��ޤ#�Z/�+IP����� S�t#-x����tɟ"�+s<��a�����Y4M@��ZH�Cv���He�N��G�"e�.���A,�N�&tyDij���]�Ǯ�n� WM��@��ELȔ�ڄH�
7V@?w���q�$N(M4M?�qn������>r���	��4�[` O�Z�	^-��PQKh��@�@!��������q��?�� ��+W?V��y�)��k_i2������K[��'W��x��F��� ���\��m���f�#����PP�N��FH
`wh���S�,*�#
1�
S��))9�A�����:K;��ii�a嘩y�L3���@����$���gx��1�k�}���6&���Iv;�.M�/���SD��3�I[�f�H����6�o9��#�h�S�.�y��~!c�)�т�]�m���_��9i�m�zC>���E�8��z^�4HĪ;�	׏��bN)3y,+��PR O�����g<>�H8�Hو�b~�R����X���tex��;�n�S�ˏ%�����t�/0c�2L���K�>߸$`���a� U�ّ��������*dYF����V~��X�wm��q&�C�[\��Vٵ����V$a���в��Db�2K�c�����/ ~��%t@�Pw��Q~z0���;������Lr�^�E��mLg�f�u6�\��,Id	��J)��^�FҶ��=���CCZ��kjkwZ��?H�Cj�yk X������}{=�o�7���u#�e93Fu^
8-Ö\O1�#M3�Ѿ͈z:����<����A�B�#��K��R�i.��\��K�P�4�����,yr����6���xgsev<�g	�Eԟ�u����~`r���~�/"�IL	�i� � ��wv՚/�]��Rq-h�%�Q��Y)�F� �qL�{j?�iw��^��ǥR_���5>9��5>>��ӧo���魁dYXX��u�X��CWW����c�	~�ǅ����~�]ƈu+�k����\�L-�>F�BUHB���d3�5��^|�-Xpf���NX˱�zp�}�˗��� !ʍnV�_9�4:��ԁ�O�����0!��"m)�9Ŗ�����r��� P�F^�e&/oH*�R�aݣE��p_X3yO��mĨz�n8͸?Ö��z����ܾ�Kw�o~z��x�a ��=T.o�$vT.Z�^b��L�փ/0�a5�Q�\/��0t.R�[}�T
�w��mx1���G&�}vC�c��ѹ^��^��sx}N��D���''?��)i��^o�+8��ڤv(�q+�z����. ��w��ba�c�=;xC� ��X�sm^h7�׷��
o:`N7�*�t����2_�"i�G�3������Nv��F�·��&�C�<������ ��,��I�B�d]���~�^XXx���Jf�EV����H}|nxU�5on�h�^�X��]Stz�,�I�G&��;	T&ofk
�"~I�,y���ϫ�Ϥ$쟹7"�m��q8��2�qv��L	n۞Z+�� I)��`˫M�Vk��(0و���;i�SY��M��/�����fw�b	��L(���O �U444ԏ�"�e?^yJO���� �T$��		sG���3�.�r�_����7�>r�·!���G8�q������� A�%p�����U�"�H(��ԓ)A�@�V�����vJE��tV��Fy�.o�b)soD���M�T�V�z[���A�h�l�>c�e�	���?�>��n9�u�X����Ν
ݕ�@֥�_{��@}�6��?�Q�EN9~����y^����l|��Y��Bskk'��6�'�O��5������%W��=���B�=��-�fC�m�9���ٷkut����ͻ���s�m@��z�ʂϩ	b����Jns�Ą�R5����V���6;�'�;~w�����4��O�(�D�J|iu��eW>�����1s`nM�'�c��j��@�	����̯յ���`%�:%�a�n���I�R�� H�����Ysh��$S]��]���(C��L��������jS��7��{Om�,�(V�˸%8HX��Į�$h��%%#���55�Vf"ne��X)��I	�ʋ���ԑ ����~�0�����8�v_'R!:�z�P� 2eRZĝT�,A��F�B�c���/Q-��GB5��v��+S�2�g�S2O�E�c�Q�UV��t>Ki�<��j[�"�%�~K�'��l7��HiNX��IUد�_�i��C-��h	j=b&�����C���������h;�)����<'�sI�l��{�c�TipiZ2�@3N�i�>���%�y�c�P穻1\������J��U�i~><?x�k�-�3N6�a������^�� S7��S������{��2�i�
��=�~�њ�ll���I.�������wO�A�À�p��i|�pJ[��\�;Z�o�3�Բn��������V��=��[�V�۽�{���p�Nh��K	Q�R�?5U���d�B�%"�.+��]�@�55���ٙ����K���FH���~�U/�d�_�k����	�N)�>f�$�9<�l�@��`�t���c1�1��9C�=�F��ۉ1�\�*�]�hᇣ�ʮO��EB)Ì]�FQ�	�#�����d�rFP#B:��݆�+YJ��Z��I��C�	NUh�v_�hni)	63����zDn�V7��s�����'S�#���%J����Ce�K�����+�f�,������\� ^KP���\}��+�ʫ�� '��Y�݅ c�p Y��z��Wv��X�_�ɭ��Rk��@"�t�;��2*��P�����0?C��-Q�d�%?�"�;��.np���eY�-�7W�#�ȯ!�K_���AP��vCo
�d���Q��S�'�Ïq�� <����P��k⺕�G���gXҋ%Yμ �3��Yo��ô��1�jưN�+?��Vc�
̃>�P='pLLZٶ���,����U��-E��MH���RL�
�3���O�w#k컙�NшW���z_�yIT���#^?�jp<�=������&���ڨ��>|����O���6�����9"~����[>b'�'s2�&��5��j��p�P@�\C�m�j��hћ���A��vtG��jy1Ǵ�W�|���MK0D�$��'�LM������x�cOnڭ�j��sM�V�/3'�_��!��%<!�
�%3��"�	��5�*h�D�P�����D�]�l��e�}�"�d��D���w\��bcdeY��.}�.<ٛo�}�u,�V"���䊑8FN�+�B�i������Q���.kDP���D���r�n����2�Y���4x�[��)��Z������|A�VIZ��m��| ��e|O���5�~H��N��;��i�
���qWk��.�=�3o��q�o�N.6��E�'����'��)Ú�b*�т�_X��o��탱�(acB���U�6u�iݲ�>k	&ah �x���)a��ʝm�MTW!L�v�\��|Έ���U����7�9�����~�)�;��c���ؠ=����Km;�B�0�B�Aw�uO{$?��n/��M�����!vkQ�#�ģ9PT��d�D取��=ew�	~�U�VfK�Jg��:v���m��k"��� ����V����yS��A�{��@�1t�rr�`� !����H[Q�F�Q��1�Oԋb2��הP\�����Ge�&��B)�`���,�/l0��۰�����b�N�{�o11�1�M���d�A{1�&6�p<��A��Ay*Jg6`���'��;r+��74��ż����p�
��˩p&�TT��A�r5�?�r=���x	�链��G�Q�h�$܂���M�E>��͹M �9]�5���"���Zu&���|�H����� U�|���b���`�a_�ة5Ld�F[;,A	'{}�%_?L
���bk֍�����ٔ�:׼�#�{AX�dT�g
Ԯ�u1�A�t���P��u6{���4�7��G�-~7Yq�/�g���ZS6Te=�^�����|�:�� ��rФ#d$I���
W��őDU�.r���� �7��dz<i]�i�Rco��Yk�D՟��c��1|�z���L�]���������g)*A��!7NJ�bp��|�,R�+�X�
�ȴ�+,�Q�E�����]5�g��\^Ʌ�f�]�p�K{�%|I�j��`(�I�GM��?����j'6�}���ݣ�{���m�F�q�\OBi�v���%�:	&�=���*�*���>�p�R٘���Q���?�{\�F��*���L�!��t� �J��5,�������b��ӌ���db����"��1](�yѭ�~x���i��m��<P��|HyA��pl��� �E88�<n��4}��Q[*�ZF� �x�m|R�V��F�Wp�A�� )�&8)��Ӭ��;��_��6~,
��Qf�nR��/�w�uf���h�=|�9�~I�p"l��Y#����Wy�3�M��{F2V�4�အ&�]rӏ�	vC?��H%�,E'J�������E0FH�-�K��L�n��Q[	7�a�~(�Mr0������g`~2�*���,=.V�tqPHm~�L$�wI*=��ϗ
o4�W�Y������xi�JX��|l?	���Hb�WY��u��Vۘ!ya�2֠�ˏ�S��ٝ�+�v�� 6�Q����~2*��w^⫙���K߿�/}K�ձ����1<�U4�>r��z��t��Drl�EoD�T=�[p�����{�E�xd}5Q��}3C��+g*at�))�T����B�V+&\WW���:H@@E�-Ѷ�@@¯C/WkZ��n�?��%lni��f^p(�/��}5P��_K3� �M��'�M�T�	:�b#�o\_��O�i�o����O�����|���($���<���z���3^z������nJ kAc/0�R���O��H�^�e�`2#k�P����YU�)����z�桤�8�Q?ҵO����-��"""�_O��|��&�i��`r��ON�h�j�f[~��J�������J������wy����mc�w���8$.��.2�g���w���/�x�mM�bW��-��0g�0\ �����8����c)�{|�{?6f�D�VU"p0"�2 �z��e��h��f�nJ��ͭU��1��\���/�׎�V��@��㍑�ff>V����I;D��:�mz���Y"h^,�,ZT)b�)��q�MP�0e��ʷ9��m� �a	���eT����B%��j��������
��
n23�0)����UzB�E�i�2���̱c���0;�:ѓ�_��ɉ��q��>�z����n^��F���[�I-A�I������><��Y��]��_�&�$�}��AT%\�o8�U���wHI�Z������@�������a͍u|ُQ��������R��Z���/i*#��L?�=e�	��)���-íz����f���鞏p��ͧu'q�q��ʒӇ�Ҋ�E �U���n������Fԅu��6+��+$a��_)��-|r�.�3����S��S+�,(�)�%��3�l����-N1�,Q��� ��v�0����0�Z�&;*?=��/?�ϼ8���\�����>^�%�~X�? P�2�V�\]�Ė�� ���ć�R�\��^�����裍���&x�x���Y��+�↪�5p�_��q�շ�O��^�J͟�����M��£}���$�����c����5���N��-rp��Ų��`0y!�	��qv?A�oa�ZX[@��Ӌ���=�Ah�5@B 7�U�_�]{b臑��p=e�ƌˑ�����1/m�CC�d[�bhD&��!�gGk��,�r/����-�l���K��,�K2�вϰ6�k�=d��B֬Ms.�_����Z��>$�`��z����G�z�H���wo��(<����w��)}��7(�հ}~̭�y T����*CD�������-77���Ɲ0�L ecqq���8�p�^�^h�TL��gq�>�Wsb�����G;uo�8R���p�ʶ����.�Y%��>Ja��b@�0�'�ZZ���%ݻ���G.l�|z���G�6nB��S��.��Sl��J�1��8���-�G��b��;>?_�{�_f��>p�3���ngg��ޭ�ǜwm��,�e}p}�`&o������{�:�����2���g�c�����T, �f��pr���z��3~gU��+�D_��3�����kD&9�(�(��]��D8�_{Z���#��^JB�è��]*�+u�k5 +����%�t�_i�do3���@H�2�1�^7���@6�J��r��g�J��	�>����#�?�H��P/�U�)�u�!���U�mR�Jm<�
4Q�94�)��@:~��XH�6A����.����U�PؑP�24�ty�<b(��#{� x68����v����0�����#j�σI�Pn5�*��c�ʳcϲPFE~|z��%r�.b�+�gμ��	~�D$�?�M2#���ꂟ>��'��o) m����h����Jb��2�Č;�s?�����f���&��1,�����B�6(㡎Lx2�XT������s�c��3��K� �! �e��Ӑ������7x�~��?9����e��מG�aW,�>�؞�"����H�dtyh��� y/�0�?�{� ��x�y[�1�?,h+##�<�����ǵ��k��ƽ�_E�?Y��Mh�w��q)�4h�O/�g��m/�0B|>!�G �5&�l4g쑖������1p�|7�?p#'� �ӏ�g��(��	ij/g�<���vN��9ަ�x��;����Bf;�p���p+�atC����A�`H�0�{b��3).2�����]qc���Ƒ��9զ���<�G�=�𫙁uk�� �����̸�����Ji$��j�#y
���u�y���&��tyެ�!�2I; e��7m]g��6tNm�S��ws��qfv�����\�S&xck�"A��8��7�yѮ1���-�w�@h4F���U�/K0��]�����%�R���h�_����YYm=����@܄^ �~�s��~����b\F��jCt�W�	ذ��؇Dr�xm�X7���[�	d$,��Q��4`�1&��N`!Bi��/����#g���d�ߒg�B��r:,}zK-�
fvvV��	��g�L�=�:�)Ŋ�t�ބ���:��JJE��A@!�,?�nN�o0�A<8��=Ch�8��WXV����0WMF<�\}���G�~na%諼c���gD;i��-&��O���SUD<�����&��FqǢ_�E��=Gr~�t@�'����U+333�bz���ݿ�5��Q}��Zf�S���u�hE��z�_�q�O=�k�8kflx����Y��h+�ze	4�z����1(�FK7�>��2y]�,�+������Ң�+%��|%'4iX9���^�9��dVk�&�M�A��8�0��x����>�1�z���*��r!p���|q�A���y= �1�ͭ�~䮶��6hVO�c0���bO ���Iyq�sey���9niEn�Uй�_'PG��bzzz�lm�,,-�����(��c�s�.����*�l'�B��7���㋙�CBK;+��X��Q nh�����ϖ��-}8000�؇���鱝RE�:���p�<��f���SYw�3�=g�wӦmé]���J٨���r#w�Э�U	�{��@q["��Z)�VQp�(���]��m��&�ʸ�5W���qx�+槻V��X؈<�+��v-G(�@R�]JWgs L�T�o3�N����t�j�򽲑�1vMMͶ�**xv�ӷ������ނ�}�{m�T!I+ \�q��'S��v��@_	��Wc�}�~�J0�. �@ӛ�#��s�zK�� H7�c݊r��C��}�2�-َ+/�HI\4bG;��r'�T�1=5�-�MI*@��du����kWJ�v�T��i�wL?���x�v)���(H O�B<�H2�b��uv�a`[����lZ��y����3{$�u�X��Ec�Mk��s�2�ʔseFn��E%%*����O4�*����[u�� �鍃��s��Q��@z�`rc�N�c=3� c8���e� ���l#
���Zv ��f�<Vqke���S�0��cZ�;V2���;ٙ�=�_h9�o�����aQю����)��><��� ��==��0+6*v����AS�(�7�s ��n���sT���y���Ԭv���ΰ���8Kj�����k� I�mlBdť�ed�	�)��e$b��9�CY�W��ĺ�3Իot�{��>�RD��`J������1������6��A�2R�j�r�-ϗ$��Rr4)����+iqhz�&eQt{������+��C����ذvuՓ)~ɽ�QJ����4s����׶r#���*�X"�؉��q�O�r߂��A����$�^�����f������]Bw��]$r����2��#��Kf���佊�����-Md���j�5zz{��w��N�04��lG�m�����<^Ĉ}����6嘲�+Ӑ��3�Y��s�n�W�=I���$���J�SYYYw���A�NLL|��rbF��T�e�/�`g��-^�����K�t��d��|�>[�U�]Up ��Aɇ$�M�p'����S�W7/�ol����@F��}���f��-nj�Bt�+�R�l]�4mҚ�����G?�ƻ[���k @?��o��#M�Ρ�5�� �S}7Kp��ҿ�u����g��={������i2�=f'+�������
���@^�de�:W�����C	Չ�YNg�`w��Q�
��S��Л�����t����m��7�GZe�l�rG�������p�6b*C?ߘ���#\J�捼��\0k�3���o�9�wT7.����#"�Ϲ�'�ۓ㶮\iF⑬p�2��%|V���t�_f<���&�\H\\�`������k�˱
���|��ӯ+�����*�� \���Q�c}�d\
��UjY#�cW���)`w3w���d�W�
-�ܱ��2����|2F��p�{䈎������r��ڈe��~sh�]]e]�s[�;�ٞ�&xXx43󱰰x�9qO�XN���[+M��!�zc�Y���~a�º�������U򴢩n��*�ܡ�W�{*C�q[�M-'�Wk�����f+�h�������BD�\wZ^]����mϹ�/'=Mb:C��d���N�5Y6��a��!���Vxjw#̓b6�,�����P4�3���6#�3�ë��;u�<�)�׭o�>�����#:��,e`m
�l����Q@?�:���PD�B���M���K��P�'}�J�v
Xm���(aU(�Tч���K��g�V�$�T,�<� �K��v�����k�煵	g�[������O�B0������ǧ+���pnF�x���N���g~R�����Ή�
+����r9f�1]�Z�Ⱥൖ^`���'�p�>��H:�"�����z��b�̜��?H-LN=>�|�7��l~oFs�)rכ~�~��R��҄�S�1�w���� )���p"��&b�ҿ��a���Av���GH J��;�t�Z�k��ҏ���c�����<e3Et�ݡ�G�aΈ����ܼ<	�iYI��4��y@!��e�FI�Tݘc���hl�~��ո��F���̵'� �^�>��9$H���ؚ��u�g9��hUk[S�g��`�bii9"�,U��o,k��t^�{�����ܖ����/_ݠ�&�h1���B���P��4��vu���?�e4��C!��9�S�7���o`�.[�����$�m�4���p�YZ~�j<���g��6�w	�QXQq�H$��ɗ�����C�pՉ�0��_��^#��K?̌f;�}H�̬�ܙ�"�D��{������?�;��y��K���Ӝ+�W_p0枘+����J+�ǒ�wHზL4F�6k�>�P��,��$Q/�70n�_.:����i��ʚ�I��k��DYfv�=e��[�P3�Hm�G"�}l����FwƧ�da��P�[��!ϖ?�
���al�;���'oØξ��Uqk��j��}!Z�Pw��d͛ر��yu��I��k����2�PY�7��3(�5��'26~�{�������f�J��S!���,F����\�;^�HgM��'	1�9!�Q̏�ά���r��Ђy�Л�y��}�� ?��:X��(߿�P��!��
�� �G��20���ݣ��[��X�#w��L��M�ѿf�w`N�E�+�*T ����^}���we
����Y����b�Dȋt ZW;04� ڏ�F"�w �)))�G9O��o�E��^�-��R��6��d7�<YX����l��mǍ�m[��� ��.R��YE�,�'��75�\�ӧ�s�9����/�SQ�E�v̈́NG����ר���vJ|�?�\����7�o`LZ��JfS;��Ō=A8QL�Zz����D ���v�|zwPP����⨄��݃����9��i8�!ur�F��a=^�)�Ӵ�q�&�Ҿ��:9[o���P�6��6�t�{)���1������}3[<Pص�ʧ�[�x> �4g �y�����A1]b	;L�T�����䦝�S($�5y���4c�yw���c�m^ʶ�P8���'v�:�n;�@���7�]���l�f=��Ǉzi��x������Vf%�|fq*�o%��-� S�&��j��W�Ŧ���'磝z����i�v���*0;,k�,��A�.���4pT�UW�(���3(=*\烁*���+r����X�;��]����P�>%a��(��4B��f��NV������'^:u��������Ϧ�G��Q��JjO �i~N�� 8L��N��@Ê?�X���ו �줾��Ք{{W�Q�4�Jm���-�.2����6��K����
�ۃ���R��*���`2',n'�� 8�t&ȞW��qM��!4aT�F"O� NP*PT{��]�O��tA��C�Q�IȑU&]�ǻs.(F$*φϓH��&ب[���� ��c${_�B�d�_��pö�AY�#��:|*�����*�g4�{���a�u^�^5�$	�_�UN��Ppʺ*�ϳ��Z�	YYc�6}��s����㢧EEJ����'w '5�1��N%gl�8�.7��\��^�ac.�s���Nmdl�#��1yv�k�R�,�?~a��|����ٵ�K8�I9�����������QG��O���%{k5. ��5q���42Bn��SL�k�pa=��s@B�ŝ�,ぺ�F"��S��=[r����ݘ�KW�âۍ_�5����NSm٤4=T�G�্qVG',�}V�5\��ʤ��M�}[V�>������Ee�Fd��@ś���!���,,��JW��w�|A�X���o_ɺ��h��XR7>��V���{zw��*'���1����jջM�@�4���|b��(���y��r�Y8'F�W����|�=�	�N��W�{��5Kƿ>S�:�(��c4�����A@�+��":�#<x�m�Ι��@�^P|��/ب{Z�W�ϤuD��q��`1頰*e�O�}�.��3n����6�qY)zږl�땝��V �W��8Qfia�q--�FE�"��=�'ىc��.K	"֬��\���g���t������3����,?�� �������?&NF�b���ɧ���l{T4�9!�U4����ňYv��V��w���%%U_�z�م|#��G�����oʝ�C�[VP�n 0���ڍ%4\�MD�n3S8����~-�ћ�ž�Mt���O���i0�z#�UbW(FR������6���_v�344�q؜��+�����*M=4Z�V�~��^3B�&3�����Ӈ�g���ư����h�7�lf��uf��[�5N�I
���}[D���Z!�V���eD�A�7إ��ׯ__K�sz��
�YM�wo����׿��?Œ�rZ�˟��-В�<e���}�ݾ��3�����6��9�)�mPrd����K
E�C���"¡�@�ݕ+�I�r(��g�ɂ},XkkI�I)�*����  �RK�G�}�8Z'T*�4|�5\�hQ"���n���IVa�Ł3p��w� y�Q�=��a\�?���ҵb���21�T���U��8�V�	Iqo[)4ʗ��G�M�+C�]�EiX3\Sz���@���X��� �P�8��{���Ւ0qXggX�ӽpaԁ���*�3�ݬbF�jwN�������E\�2uc��n\_�����U")y� �>�E\*G>��e�_�=w1j؏dt�7�C���jBH����Û#�3��Umll�;8�a�_>d��Q׃3��;�G��/s��ɚa���T��x�
K3+[ н?M�x�/���Q�'ĳ���	��O.�ؕ��d�l�oi.�k� Bs��2�X  � �zGw��1��a���E�222�'�E�����<ͥ����{��4��N~#@;��K
�!Tl�N�Y7��X"8\"�=�w.崭�)�;3�k�㝚�_^�Um��"
6`JK�ΞEG�5���G�7�m��lF�[S��Φ2ӉU����1{kz����ۭlc68iaGC7`�͙��VV��)>�ו�_�s:��]H�~���5��^���xj�Ʃ�on�����+�؉�Un'pX�P�X���F0l�K��9��CW�'N̻��a�+�S����<@ĵm���������X�o�6nx"��.�L5&.H���Ӭ�ڍH�����B�M?����kc$o���:ۄ�Dp�߽3�>)�z ���myy9��dd����D=׭̔[��(4��뻾J��}��Sj�L��6�z����0��P�����趷��<A���5ad��qL$
+/�wu?�̥
�0?�=}
|�s�{z�{�[N��f��H��x;/lA�_��(BKK��D���F��/�E�v�p�d��#s�m��?�G�@�ɵC}��Q.��?6<�h���q�vy19� V��ld0�������7��LH��,�L>p!��L���(�Z7�����:��on>M>��!��{���@Q���n&����<&y�=�����o|G+<����'rrSx�aiA� �	y�}�{��~���ڸ����Ez.9��wns1lO��� V�8gT���U�ɤ�I>��o��J����� �rj���%�Z�}4��1x��u�����5T�We�]e�%`��6��R���ٽ^�3u���sByI�f����
R>+������>C�h�$����;��`_Gե��K@��~� �Z�?�<S!5�PVs��C��<L�L��}��D��J(�&��yc�蕡x8u0H��P7�o���� �xe�k��;�W�%_'V^-~=��ޮ��JO���?�b�߉%Щ�>�d���zY˷o���!G���I3R5,ᣣ�!�PY�c�����^�|�0H�_.@zK����04�)�{fV��B��7�|�u��ņ9���Y���V�3�U� 0/f�:%^aN�
~-t#��vj�0����p�3�챞�蕊I&��w�}�s�id����R��ގG�L.����;8�F"�V&&^Z��֖��?ef�3T�Vk��Pﮰ���9Y@< ���v1���X���?K!3��"���_�9��s�<T��؄|�G�q���`����2�4o3�ח��٩��M(2�x�Ev� T#5�4t��{5����=(T_�b�������� X9�^B��k�,���]z�G�4�K��D0�r�N666�6LHH(��|�av�?������)�9!࿅@R4��SL�Eh���H^IdH���4�9s�$�Y*����F󍝨���f�;iAY��Ƞ���4�Ó����M�,r!
1���L���� �B�,�!U@YlR[�sب9�ǷyC�Zp=`�a�������y���a*F��Q<$M7�;[��״�l��%'h�$U�J	�NX�'��\,ot�C��][�Zݓ_��-4E�{�7���{O�j��r���5�|�uj�[��n��6.$�����ٿmn�AK[�썕�^*z�L0�����[OO�����]��rB�n�E��3�}-`9�7�@�l?y��)���~�L�*��������c:��!�G���_!�u�n�N\]���v���	U5���ol����y����S�I����ۀ��A�ĩº]v3����#t1�l�����LM	.�I{}�nR�����@$p�wv��u<���რ�ﱩ(��#;+�4��hR��$M�m���H
���}y<���~��T��QRvB�X���Pɒ}�2H�2ȾD�THv��o3cϒ�dC�C�L��gh;�|~��z�W��q��������}���r �������3�޽CʖًX��W�AN��s:;;��At|w������qʉ��~4�>
k����b�YE��Ƭ�}��A�C�npf8w��c����Г5U��~QY+?���16z�#Ǽ�BK/�O��D������`�Y�_汿É?g,����@�ϡ��mԵH�3�jq�	r��LJ��/�b,�V���n�/��<��ϳ�\�~�Ec��RQ(T!_�`�Z�~���%�Fs�,�	��Ew��&�Mf!z��fO_#��e8�9����6��d�)���^��Q���ƽ>0�y7��3�C��S����>z�=��g�����e��n��(߳E�,�Ѳ��aTE���b�{�"O�q�VG.b���Q�"y��A�ݢ�	l�P��i���Ǫ��o� ���4*:�umxg�v��!V�l�]:����ϧ���C>:�����J��u~�(���n���#�ޯr|A?�����Vnd�`�U���q���?.n��R�(����Nr���W������;��C�D� s��ŨtG��=�gw����k��,sF'�{	�����I�
?�뮬�I�?YT��Q�#�G)tZZZ�oI����{�[X{	���5�zF��_�&��\c�R��1�a�X[��|��1x��b���ـ?��b�@`74z�i���v<\�д�~�ՓyG�)��:�5[L����r�&��ݣ4�:k��d$b
v946c�E��oG�v&fF�C����$����A/�L����T�+��JJB)Z�tijAl�:�p;|Ȁ1	+�-Y�<��*�Ճ�8��~ݨMj��|׀:V��b@���϶Xk���.�!�LL�k.�O
|�%ͮc�P�p���rP�(|s��ͤOR�(X�RlBѭܰ�$���{����(mu��"��E�����S'.�H�m]}�DΤ�}��}���̪�ŏ�㋎�2�����������%s>q��d%���@T��LQ��cuU:d�§;DhsV<y2s��
�h�����? qn�-���S��z7!̹G�dN ��]w�$����ҿ;�'X'ł�s�ǀۭc�z)����$ժv�}��<l�?&2�����h�ǌ�VϗF�Ǡ,���z�
p�Ԯ�D]>+/R��b\��32�����"� P�"��t4�X��x�|G��a��0bR�DG'˜5�ꧡc��p��!���ޝ��/����d��Ұ����>_0�gv���-��� }���(C��ua���0%��[N1+(9%<)����M������o!�����h��r\��M�V��ɿ������H��i�n#�.�O�������j�'��Y�N�?~�%�Y��C9@�2�u͈�6%�1�;����O���w��@Xb^�v2�3e\i;��(�)�FνE�T�c����Wm>�%a�0T%[,Ձ�չ��8��dvv��<�%gFo�
�޺g�<t%�#]���0�%zB���l���w��_�2�|�wF����.Y�����ypu��Z�أ�����=�Ф0���dŢҽw��^��@��Q��]��@�?H�@�$Z6刕�zo{�#Ȇ:�Qo���?+

���Q��3~Ijۧ���p���ݹ��퓋���)"Q���v�|W˥A���dN#C�L&���y�<�4�F�����|�Ԑ�"�� ��K��G`BC� +���M$��x��C�-
�Ȯ�r[�_��;O��ko��ґg����p���P*@�z/����s�:>inq>#ձp�TĀ[��F�pV誛��'FM���8@s&��O�`QG���t�M�s��t%p���4�`)>�������&u�<����[�P����L����������8Q���:9����]�[��^���,/OELx�����hP&�s���b�x/� 1���s9tH��_#!0�{��NU9��n�����E�����A��.�� yl-�4�l��W�i;���ϵXNPT�I������l��oau�Q�Β�:�h�up��ʻ�]�su����� Iy���Q�6Bbb(܋n��M����N��ҒR���V�C�*�!_����{֎Y�<��,	2%B���fg�b�7A����.�n����XΖS��i���A�4�(vw����a8xb�a� 4c�{�$^���T�����7�}��PD1tg�<�<+6J�Jy�ϝ"N�*����oݯU|5�C��HGt���e��3�뷦�S�KnR�/�\�6���Z���GYb����G�l�AQax�� ,��(9��g)�c���t�09��@�ΧFJ]�tȆpr��`PCJ��B�& ����z�)ݐ���� �8�『��U�Y�>QIK�"k䨇�D���`�;D��T�̀s?��?��P�ҕ�K@\xD$�y��0�;YT�`ޓۼoቛ�E׫�����	�j�ES9�Կ�Έֺ�0���d��-�u RZ��ՠ�j:]vg+=���{����o���+7���:i�O��͙ P$�^0�qrr��>�����������+�$���R2f(�"���bF�ً��%�CE{��V��*i��4@�M�i!( ўޙ����6G3U;��_6x���{0�2�G"R��m�آ�O��[�od� �@^��Us��lt�*@��^����7�i��$����L��qMB%ͺ�U�3{����;�ҡ��)�|��
6Z��fN�뾠�.��Z;�>iA��UaNk��}4t���1�g����ͻV�zrR ��9 >V��]Y'c��ukB�4���i������_��~�49f|�$��4�?%gG1׺tn�05�d��th��G��V��(��6�kK�������K ��SL�9����`�	�q�uT£�B�V.JE��+��<�(�x���B��bL�Cfe�j���?��������C�=nβ��s�8�:2�L�=�D������c�P1��&=�D(��C��ɤnCڤ��;�ł����X��'�lc��ߦDƢ�c�g���VEN�o��u� ��b��e�|��{Z�O�����໵ �:�q��`;��3��kPǯ;� ��,f�܏��&hhh$��ܹ�Zf �<F9�������Jd�A�p4i~pw��n���t����E���%@�/fk*  ��%�����k�sPP��&��g�/_���ěߜ:� Ёȓh�]~���]�c�K�<�܉���BE2fc�15��氐��[�*�9#<00�G����?���V�c�9���Q��ሒ��nh��1�E�j�x躓�S*9T{CJ�������Pi�:g.���������I	ֵUYx�d�g�̭��~t��icŊ�"��cc�[6�����6�<��mmà�9�4����ǭ�nQ��o�;�'��HCC�W%;̻�޽����"��ˮ	��5b��m�lJC�т5«A�7x�gx���޽���X$�,��{�7�دnLá�[}@��ų�����S���~R���P�(��M���#|@���r���*��������cbbb}�4L3@X�U�¤&��fF`��2s�,�����[�{�A�3(�P���D���.$�@�؜�k5F÷p�����N)FO��}E��AOH�EUtVW�F�I����S'�J&�<�O>x�@n���خN^yi9TvƱ�#�F�����y#�(�,�t�{���NsjJ� J��� #�s(�CB�������yP����O����{x/��S�iy:�7Wߒ>¦ǖ�\�OT�^MM���eАpW~L2/
�Ǐvg1n�R��\�S�ʛ�yg��@�D@X��0�F3�6�֌���a�(K�x�F��3����+$#МR��;�Ec��oW��4�.�n�����S��р���i�L
c��ӧB�c����iw��1���K"X�L�qnJf�(T��WFhUo�mQ�=�)F[<X��U�ڋߙF �矪��g��������A^���� ���?`<�P�-J-��f����u�cC���|�␦� ��b�?Q��*�ߝ�4����t7�B�ҡ��C�+>l�������:k��}�Z�#��w�d��"����$�k}1,,͛�]��#`�*�`~��eVPW9�R��K��Ii�!��z���%�.���
S�0�q�w���ᏞLݎEt2�;,�?"~�(Si��k"֫O��� �� ��P؛�zbp}ee��1g---���,�� ȑ62�G�"���M�s�_F�wx�^+
�r@ �'m�W&4����j:�6M[�F�Z��񵙠�e��1�k�Ldˊ�7��@��|��꧷��.-��*�iw@�k�2!�^�W���#�j����9$����?���4TXx��h80����>��<�������0]^�	�t�8�bQ�-��������'�364�ħ��R��H�����T�cw�"+����D��N���)��� ��_ݣ��7e(�w� ު��MOƣ��>�>�[2^�M�K�'�mNh�S�>3�+�5�����,rK�֊5	�w�lo?�����c��.Rr�7��jت������ŧm����#�w��1�0a>��p����hg�f��n��FB׆z5�s]\�H�%�ƹ{�P�1dv�!r��1B�W�[+�#������|�Bקm̿��.wA+ya�nT<�6�00u��I�A��n��M%ZCi]�ܣ|8��˻�g�(Ϧ����ث��T�!at���O��,��;��.r5I]Q�7�zй�O��Z�Ф1d�ߏRٝ1W�ڦ�#Q�$-T I].?�e5P�����ԝ_d����t��c�E��,�ؗa��-*E�i�
�t���+#�:Y�r]�`�U/�!���-���HV�N�|�D	�4E��J��'7���Dt�l�rL�\Q�Xww7yW�<���(@|�iM�ם!U�H�R��f�E
�m�g�)�o���v��P.=e��;S�Ȱ�z����#A;���w�,w|����З6}HC�r���;;����r6&�$F����ɿ���Ԋ8�]H�*x.�m��+��Z��.���\���UK����M���)�ixA5��'w8�W��0U)�5X`Q��`u�v���kR�-��9��	���^�w,�Y<S�k�0�>-�
&��~�]��bsR>n��
h9@���0����=��Ԅ�X��wM�VA`���"P�6�e������[�3e�v��k/ߡ������d&�P���Kx�γ |�f\��8�p���Gɑ�oEw}����x��{�
q��~8��mwO���/�5���={*%g~2��y"�CW���ǂ"�b`���J��`�@�#C��q5��%ڨ>!�r��'�S/3�*�K�^�ǁ���gh����g�n�!,M�"�z�$�^�z=��o����xZϞ؀Dm��O�r� ԫ\��E(p�Xݳ�i��M{,������]�ef�Gt��J^���v�3k���0A?#���<1�L���x�^b�^gx�{�e�f�W�wha��MLLLuE�k�0�+�S��'B�|0JJ�,��SV��Fo�'u����t����'��p��Cj����h��{z�9}i���+��H$𑗊������F�UZ�y�M���7x���@�F�p�s�x�g����mp������KYY���y��a���TxSX��4K�#�-=����y�Ѫ~��r.s!��7�O<I� ��h��v�#��QJ�}�Zef�La$��o�P�!-�����Ҽ-uJd&sw�z_<�I��{"�?

%��J��j-�rltA-ϝT*]��ʜ�s��g��&�;�ao�v��*����.�Z�%kv�61)��S�W]
��4�C�R^�ENݕ����6'�xlc��Gj�ňC����6�[�A�KD�ܶ�	�pr_��7��*�?���?tڢ�e���kpǫ0�
A�J�HKK����T���A�Ԝ�S�}�+uc�bq[����o�>�eC��9w�������"�}�v���:#�+|,b,j#�4�/�����pJ@���vY����@װ��j�<
���й�n�Ckm�{: Mb��᤹���U��C�f��_���.1�Ș�Q�D��uA�:ޏ���y�����,��32�<���� �L'U}�gA�5�5�~�<�o����[U	��n�"� �� &3;{c�t X	Y�D:I�)ї"CƧ��O�aR���;���g�82��Y�[�~.䉤 5[���;�Y6���M{��$�?��ї�G�7��g� ��|�X�\��%��a�8zk�����#|�^��r�~����-���n~�e=�pY���?LN�~/#r����*K��k�AE�|��r�Z�|rO(��W3M����HH�@��6L[������ّe"'de��vk\YUl��I������ҧExsI9�QO"�pO �G ������2�{�ǖ&N�T�km�$���.�U�D�9��_�e�r���b��iA)G2ijf�k��I��'o_���" =�?��(X�jߌ+��
��+�����`���"���G�K���n����ν��y�6'0X`hD'\+��#4�	ss��cK����m��q[xf�"7%~��c�l��1~��Z�<�����\L�\�$�;d)��}�
��@����M��5���Ռ-�񢬹Z��mZ��fm������y�;�#��5'�T�*����1v��}��}�a=%���O�X��uA1�]��o���U��Ax������5l�۔�PS���SV�v����)bV,���[O(�ۯ^\�XX���]�0��ÄR*��Z���L�&���ϴ^2��u9hf[�m6��X��լ5��p�bU��,M�:�lЛ�b�<p4�w��؋��pzG*��	󈹗�+�9��/� �"����N٠��&Kq�tޥEϳ��0�ط�w��t�+���V�#?�����=�L��I�ܞ4X�tw�	f`���s��W�7�PL�ιb\��
���8�u1�Ht�ֺ@I��Q�۠0꩎�?� L0��J̨���3Z�J�����?�-�7|[�$M?�#��p����L�ߋa�߇j��0���'�-�l�j����U}��U���PO%���k|�͑�-����Dq�¦!_X$Q�{�,�����9�y6�M���S�H��!¥t%���B�^>�",q�>ece�x��"s����Z�a�??w6)h�e}���1������~���˒�.�ΦQ�C���"�!Y�-��Ds��N4����F�)g�E�AMoqJO��z�Ȟ�W�F���a q
��;mVo��^T�����g[z[^x�|M�
��F@�"���%����sq/�`�d��a,��<�[�������b���ĺ�6럛�.���O������:@[��m-n��v������-��0xj6����x�a�^>\��� ,������&�V����0�����j���7�.�~����20.=D�:�+ݲa�_�!O
0X�� �$6�[��!���!���ke5~AueI�&�aW\�e�.َ��y����wY�0ib�� Xu���`�7��t�
���PP& �o?!79t�\9L�aU7����~,��sv����OhC5��&�s9y� Gh������"8eĞ}H-��&%���E1�5zX��EƦ��#�Z
�a��K8��*ye��ޢk����Mk��L-w��K��v�'} �"�&o�TM�����@`���8�|F	E�"g�QoRCٴ'Zvf�b�8�d��<��5z�=�އ�0Xpx�X����\�G�h
'��N�	�D��{Q����c0n��郓T
��������~���|w�b`4t����g�FD5�#��E�`�!E㫌|ma�<qD�t�-��+�+�����ŋM�-F3�3�ݮ:��=r�Cz�deWin�d�Og�g���6��s>��9כ�﯌b��ƫ> I���,��Op��m���j�^=9�8���I���˶_/Ea����E�e���c ���)�ŝ����tZs�ƸE�#�P�Jj�2�;Yzf�6�9�r2h����̫��<{���鸻(��X�+�����b�؜ļs
Ǯ^�aggGh�!���Z��_�RE �|y�m�@񛫆iX�X�&���ڠ����}I�7k�K�����v=�y�U"�|��Y5 ˫��R����)������^1��]�9�h���.x�w��Ä�m3�N�R�.�Î^��ԣ�w�-��ڝU�%��&:���-�g��W����D�P����ii(�1�g�@q�d��e�9M65�T�-9d���1�G�������g.<�Z�
C�w����k'U��͋���8_F��Ħ�At�@rw�=j��y"�<����D@���*h:�r_��/�ʂD�
�4�M*�������&X/9|)���3�W��?�k�9H�fӸ�,}��A�"�omu�D)�%��[h�#��(�`���I�R�Rk�<b���^�h�K��J�r�/��5�e-hǚ� �~#]��d��{:�u����r�ڃ�R�4�8L��5!�H�C���mm˾mP�	��������ך�9b:Os���木�FᴆA@���4�փf����D�:����qDTi�^k��}h�P�rr��l�39S-�!�~�~s�*�b>��B��iu��w�(�2q��O�Wr�0x��ފGxޟ�(#,���!DA��ȑ#��}��WJp4�xk�K�c�1��L�$����[��-��t8�v5��+M�U�ܿ��9�\�����A���,�`GlvOyp>Q��ӱ��K2����H��'Vx����SՐg�F�h�bx=���P43�'�,�>&��+5�Y<2M99r��K�O�=-���^���&T�l��p��} r�����ϻd�X4`�P��G�&8��ŕN�nI�u�6X��`�!�a��ee�[��l:(�OےrQ�y��%P�βbxv�Ma���+l.��k9?�f�ʎ�qAtׁ-�I����	��F���[�T���3�;�W"�����O�T YJnm��i���̴�k4��i��7a���%�o޼���,! ���w��XI��Wp3�j|7C���-?���)�z+N�}�]֘��[�&j�=`��8p�������e�h� ��
P"�?�7��V�����9��-�C{�P[E�u<>�G����7q��<����fI��?��߶�< ��>�/�)M��[�pڲ]�3�uC�D�SL�6I�_�˱G�Mm� `a����;x��d��"��%��@(82�*���^��"^�(,����n��6���6��d\�!�O��R�NV�c�k�o�?����]��~[��-\���yD�Nn}ii�Z,Ǒ�>fM��эS�jJ�9Zƴ��khLEiSJ���_�P[�R2��S��ԍ%��$ ���*����ˎ��։�b���� �u���'� �ih)����u���)o�s!x�N�R�v���
|���bKD8��z-�ڰ�#XN�?�v���F�d[�2�"�Ḣ����ї��1Iͭm*{��3 O|�Gd����Vݯ���;L�(��}Z&������QU��0��f@�+	�&����:�]/5_9s��);�gf<҃?�^� ��K�Ozc�L/�� �Hp;Tט�/3l59��O;�x����tt�Z��9�)�{4R�d1Z��64�� i�d��R|������x
O�,	=�6^%W�<m��H~#���Om��z8�D�w���s��TO�� �S���%�RX wAtQ��b����_�e�����$��4=��{�S-��g���)�ߺ�3��Y���Q���dJ5ݝ\��Z�8+��Au��0a *��u)7
�N����5�_f�G�m9*��ӁH�^�r�ޑ�M���5s����!�?:PHQ��pe�b7�t�`}���]8���5B�{��d,0(o\@1�����C4�ƬV���a
�xRW�*{���~5�8���/rި�CC<>7�h�	Bx���.�<TC�^����Re�<�5�j���M����:`xj���LY�T�\����,�6
��e� �Y��ެЗm��<�I!�`�a;�t]:����O#��EcŖ��=������9F(9��O�>�tg��,�?��̊*d)Yc�I�m3�#�B�)�mY�[�/��^�2�Ґ`�ѝ����#2#CԽ�RŸZ�+�Y�=J�J�����������=�0<%.{r����h��D8�s>]>f4� uU*�Y��{��ͫ����f ���(s�(��OG8X��10��pR�����.^U�E+�S�<F�Lu��mi@�x��[w�=�e���c`a��������}@3�=N��S�>ٔ�P�T�e{,��r�~��3�-�L0��r�⩏s_�(51t�����gG�����A���}���x�W�[8��>t�]v�4�
gӤ=�P����\Tv��[���F���o��k�2�ܒ������q�� ���#\�I�]�����S��a���nW�R�rZ��};�-�K�����;������u"LMMI����Hl��:YE�^��*��D�Â̠=����zY����c��:`��`�=CM����=����}���[���[ Al�6h��7�4���*�K���~v�hu�����8�����_��K������a��no4�,��u|��!���w�:B�M}��-q���1���)f@�;�I9�4F�w{���)�D��Tǃ�k�j��}�n4!�Z��(7>�����-c���?��/^��Z���\����;aEnA:�H;nvP~J*ϙ�zG����M!�s�F ��C���B�i�5.gB������|�
�4��
\Y�Wtnbȧ)[6�����n����x�j�B(<�ܨ{�(������,.���Œ�H���u��%{ M�����{�}p;�2+��^4S��Q�RB[f��k�����uCDd�����|kg���i��R*C���ĥc�Ӭ�v�Tn����Vs���tćq�1/�v��o�\� �G/��Q'�"'�U�JI�I��Yp$��@ũ�ϒ����p[���L��g�;
���j��E�1L;���>i�{[^����(=�\s�V�Fʹa�te�������$s�-)nA�!K�0�S����z�c��7EK'O�*]v�����k�9��~ô^W�c*��0��n?�k�mݻ	�Q�X�|�е����a�=*��_ؔ'�l�:���)�Ya�!6�ẎI�G;	�K񦙼wT&�n{>F]�����1��`���GQx�q�0Q�|5}+G[Nŝ�>�T��-�~6�LX�ሃU�,Ο8�CK=x�y������Z�׏.էxh���ٲ|@T��8���1�����Nɡ���h��Z�Uߖd֛�X����@۩�5�fj�oa��J<��E�Ueg�UA�{-�����D<tbf[(6z�U�9�_`�J��}w�6+��gM��s�x�Ud&���s�^Q4�x
7Ie��1�����'Þw�9ȶ��l���Y�=mp�������-S��*�y�[E�hg��@�	�a�\�غ��V7�v;m�v3��F`��\��[�[� ��*������~��*�4�s>1��~;����{�ԇ_K�����g?p��4�<9f^?SY �9�iB^e���M�ɢ��Y��J�Ɇ�^�ǂ��^{T�.K������K�ÉgH��*�$/�_n�΍^��K�CO�Ҁt����ة�ŋ+�	�pB��&���e��H������+م֭��0)�V�R�:Ä3���Z:��|��:���ܳ�����ϯ�0�o��Z���πtCI��b���T����[��9F6=(���D�6j6G#ßv�_���3pDvZ��ʭV,��]�I2�A'\��w+�y���Xo��i\X�i��B�c`����z����a7B���
��K�/�ZEX�!g��}��/�-���	J�ǆ[���'���5�3���ڣ.x,y-�RxR0�Y������>��"dJ�.mG���OӬn�2�>��+?�Q~���!ϖ?��ޤ��pq�kɫ�L�����'��ˤ9 �M� �u�<"�}��,Ƥ.z��U֗{Y·���68����1��Wn;�����x-�W��^�E|x.s��2��P��0A �?^���i�a_��LV=w�co�]�O[��WQz}DN�߬���!)�
�83�8ݓ��U����:Ḧ��XK1�:M'��~�����C7Z1t��FaԻV}Y+C��0�H)�yf���w�0�rY�c)�[�-fs'�W�Z���
\���b����#�4�D�B���rV�=1�u��Պ���y���q�Z����FQ����]������Ē�|aW���'b�;�ε����n潨*`\��AQj��|�/�9F� ���6n����@(L�RV�_�v(]35�8�+G"Vea���0�g��Qzb�x%�+����	��Z�$�$3�h�,⇬D��-����c��F�_�R�dN��GI>���+�8��P�e�^���խ`O���m��u Fs��c�vr5�K�=��_��z&��?*�W2q:�����O���\�j�^l�2$�|�p� @�Kd }�a�uO�_�%�tu�=c���'��4C���-��ִ쫥���^��g��"�������P�P�w��i�����6�w�Z����uB�@eu�#H*ڨ�N� �5���$&�`����X��·�+9�� ���^N�/Zr �>ճ�W��e!t|\hV�o{3�K������.��)�8�sgp��<����+mz
B�`|����a����)��h4���-�<�S��:�B#�����Q&PqE\���OV�IH#�����G��6ؼox�-�����߉�[����s�h> ?�4�����}��<�N��E��K��e��{V*����j!n��.-�m���Ɓl��e�Վr�@�Ig@����zN7�a�&E�L���Oې��SU�M	�\�މ<����E?��|D|�~��E+ˤ}�O^�YF��b�ٜX�׌��{5;��D3�W��"�#u\�mQ�����U���Hq�Ӹ~��1IT#];���p�t>Ȍy�����E5�&#l$��ֹ� ŗ*MPe���ȝ���6�(H!��&�*ث�4��!&�U0[�g��9���5��X�@�G��6�ٯ�b�_˯��w�^	V\Ȩ7����q�.�(��)$�^m�5��mpv+�:�f%�1�0�@��֟�5^������/zr�ԁ¹�S��rV�0�3�.K����g� m��.����f�=X0OT��;r�������iJ�31\�azB:��"���:-ԟ����Ҧ�kEv�X������9]�&?����ΑZ4���a,H4_c�\�O���y�s2��^!��WU���Q3�^v�.n ��"���7W��3�݀��e)��!o���Ǐᡇ�dw����hh�d�JN&�>�*=��U�(w��H�n����9Ps&0�W	��Ԥ~�'�tO���MQ���i�Oظ��w�,`�Ä7�%8���0��Z!�S�r��\sj5�P�|���K󈰹C�O\/����,Y��kՎ��.ǽ<4�xFx�LB�/�m�7�Ƹ퀬�?��ӵƳ�J;]��.����㨁���c��wӐ�d �/��n��v�:j��NZ8�����Wn�0;��/���B��C�]����S��f��F�̞�`M��O��tB
����6C^�]���'��ӽ#ѐp	D��KҾ�������`�z�dNhk���hX��R"t/C��"�tR%�Gp�T]Z+L��8�h�*m51��7����y⍬&�}��%L��'�?CF>�6{Ϟ�(C�m8�I��s��C�Ţ�Ů/oE� �� �r��LZ�,�۪@�;sd�d V̮E�<�z�"����C�m��H���®���۶V�+��
�F��\���3��o�܉~Q�GC��<��(�W��v��I����wfھ���ȍ�F˻oH@��Zg=GvG�<v�0��+�o�߿-߷'���.c�AZ��\F̿�;3ҕ"�rQ�s)�;���-eΒs�-���,���y�09��
�ݢ���
��W*9>0��>��m3L�#����.UA�8N�_le���}k�C����1(���jω**���8�������J?ޓ�Y�u��S���._X'�\p�q\�)D��8O�'�t�]���JߜMGegPέ�T�'�Q�d��������s�w��hd�ү
��1K���bW�,���ǅ
 J�q��X�����K
���^#�A<��P���mߋ��6��	�ë��1�������.M��HQ�f��G��f~�W�+3�H����1�bEk,��kT�=��T�!�T��7;�,Q��ˌG�������y���s��\A�i���5����3���3~�r?� -k����ǣN���ŋ�.�8���Υ�9�����|Y�� �t|�6=�pI�Ə�=?F7׊~���t�/�����ç��Ķxī$L�ē�t>	[+k�%��C�A�����c�р��@��,7�I�8�YY�,v��*�U(�5==M�}�0X���.�i�.�o�Ci��r{�Bn� S�d�E,�	�T�jt�x�I�!ː��I���d;/�	 �� �f�ޢ yc5���9!z��L�?ە���D�*�a]o���.�aqPt����>��Ƨk���:�J"wX��3���i�\'}|v���?@����*y�נ�����Vj�P���?�G���ȧD�3S*�uEQ���r\Y@�ʕ� �k��ʛS��_c���C'$$\�x�",�(�� gĆ�8�0��yWcRg%\�D�+��?͌(=l��F_��g���J�H�n>N��P���+̿���Zv���8�e)���A�]P1 nV;�9�c͌��9��1�S�*Q^�!��dJq�'�DV�Xn�o�C�U�" �E�����O^��l��ê�{���kR��5��E�M�N�����9��\��C��P�P������u�68i����y�؜��{�K�?U��Nײx���Z���3�h0����~��B&"�H�-�Q����;�}z���E�I(����[� ����~l.������k3��B���{ ���
֞`�S
'��c���8�z����wp���
>�:����
����}�ǉ����-�����7�u�8(�=y���M���A�yk�"�j�Kpe,���1�&�$Oa�e�^̦z3��F�s��?s��ÆH��R���)u�R���o��q��o��o����ףՠ�	^O�A'R�a�B8���=�'�lRtGQ�,�C_Z�B��>a�Y�����9�;��Sr�F�.ߑ�����e�I�﷗?la1��.�r���|��ڄYl	
��B�P��\��X�j/�z�(�Iy ���'�k܈��;��
C#�ɒZo���@������M�	�~�@�n<7GK<Y�\�>qk�c�M�f9�g��5�8�,��ߔ�?��J�Pl�k���~İq�A�]=O����<d�O�(�y�L�y����^^���lz�?X�ޞ,H��]���o~���'GL��-�Оp��m�)!��й��;���B�h1Y�q�sȕ�5���?zV����WT��	�0�\9����<�>u�<����bP�*F�J���D�� ��!��*����a+����A���gXax�[��o36A�,۠	9�Y�Fw��F���q�v�erj�4ʉ�V�EhP�����z��+������Q� ���뉻��n��j�DXs�#Zio*�4ꭝ,G �W���/���5���澂�4mf]9���졘��?�d5lq�MP�jL�>��]N_.K�p�*fcP������ ��f���e�`����Im�I7v��?���Ak���^��`}����jx�2��	�i�~�-(�i�㇂d��V�0���ɓ7���_���Em�u�|��^�`#��i:y�=���GϚv�&z$Y��Lh<g�H֨I;�6����З	�F"dYl+py1~�Jl�ϔƟ'�v�?4�*�d��3:���$������M�"-B1z�賋T;��3�J��@�ɶ��ji���w{�TM�#^`C覚��^&o�兟Y�m�����β`��l?��$p��+���]S����ۣ/^d�H�rdEw�m��Sür4;q��n5��FK� )�θ]]�|�[jȋʔ���'��4��C[��o�_�$�i�)���h�z�lD�G�~��:ǬKq4����m���|���Kb]M�M���}w�r���S�⽀�.u���2`���Y[���Wy���$8Z=﵏��L]$W�x�_Q�����UH�i5g�:������>�ek ����9����y���=��74�0<T�N�/ ^)�-g֛tI��ҽf�|���njX\?�����'���{�z�O���B�},�v���_�.Ƞ}��'�"/�>��	��E���x��6���U`��Kd�"��2Y�c	��X���)cl��$;�������J?��'����yL��� 3��S�^F���ɛH;����Cr��?НX@��~2�&Dd�˫/'II)�9�d�����H2H=�V��ىX����]��?�m��<ˑ���/�F(�\�m�@�ҍ&�Vr�<��EA0��տm����w�E���N�~�t�Y��C�m�����r��oB��`��NjB�$ڮ���;��Z��+���ǹ��v\�0��f�vod���X/����$����e*�����bh3�}�ֶ���W� |ܮ&Lr����m�q7�B�2�`��wܫ�g��ٱ�2\s*�w�������R�G�+b�N�?���.�n�����7��R\|[�v/R�?o�O$�>�g�Sԏ:\�ڧ<vܫ�C�"�w
z�iA�w�.1~����ՉP���V�)�IWv�Dad�{Y*CnD�yl�kY�*5��zJ`��> @�B��^�@9l5T,�PPF����t%��բ�O��t%c���)��Q�V�D'u�!Xmv�F��>�A�<�N�VˢN f�b�z�o�V!ϟ��ǘ�R������(��ݣ�ޙ�z�r�h�U���C���Χ��:n$�
WR�(����.m�_-�
(�� ��P5u�;������<��t��x�2��˼m�Yk��W��̭O�.o��nvM��N��a�&/G(�U��eG[�\� j-M�Hu?6Te�D�տM����D |u��A�Q�����ja����_��X�r�e�V��_���֢黜948��7�S�7�X�x�nz5��V:�:d/MWC̅<�-@��o�wx;�xa(��>���X����#��@oD�}����O�I�5[��e�������gSM��j�T�(���%�n�`Hd�t�.��d[����EyV���7��8�T4����/��O�����: ����1b[���k����mS����e�.�6x�[�@�za��>(�z&$Ui~�H����0C�0����)�Y�����$D�����6W���q���Ygl����q��^���RZt/2�@F@�&�-�F��}Sw��1�#c/H �=F<�)�A�Ğmv?�h!�;�N�r �{�!g�O0q�g2����Oɘ�B>}?-�-z"2Dh��I�,;���3X�ǜM��l�L^��!���Q$���^}��q��1Ņmp�r��жSj�D�8�������8�L�'W�k_�ކݦ-B�Y"{ٲ�D��k���L%�)�Q���,	Y�P�}H1���J���<��}���9�9�9��|��������{wq�	�K�{1cq��tWг�nV����_���u�4NOu;m�U�{3�	���]P����a�%�_������+���{��L��M����������q�� 1A;{�Ϝk�3��7�`X�ђ��ݠ�C{���R˱��������5 �S�r,��1/
"��t��S�X�v���X~�!m��1��mEڵ��(����|����[n�B�k��'�!���,e`9iy�a��?d�??�Uoo��!t͆xR��{�|��]\D�Bc9��ͷ/�0���L��.Ž���O���Q��G/YR�C������*�x��?�(!�$�"l���D���JJy�t-=G��kC�w��g�����k����X�.dGX�_M�ɐ��	�	������1A����/	�k1�:��R@�C��p��N(��i+�<�Q����ϵ�z�`͓$��2��P����f��c9h19�]2b}}���/��׿J}��m�·2]�[�$Jp��)�$��?T�8R�xɦ�h��Ќ��6���o3�T܌���(K`�kX��B梓sq{cY�������>���恋.���@��f�J�2?V�Tz�D~�1�]�!�;xrcDWX~��<�A��=@j��٢qx'��>��k�l i�0G��B�f��J�w��\�,�¥}��rz�q&�~��dG�%Q�M�Ɉ�-G��g��p�\�:� rN����d ���v��6��ũȋ�do�h�hF�9N�ty8���tퟒ���F7*�̵�D�1[_'���tiyP�%�r3M-�����Z
}�w��T�Ny���ߵuD�%���y~'`��Vq�^c�W�R(>P����R.݀,��W;zk�Q۱Ih{T�R�z[X*�V �@�)�~����#��^�=���Wnm��[?=p&�}�f�Y�Y�� .����H��V�>Eʕ���ꋲo	�O> c���fNO�g�D+�޺��y�Y&�aķ;aiȗ�ϽXn|!&/(*%e�8�fQ�)l�F��x����o
o��+B�-�U_ b) ��'&�?�t���ř=��&,��R�*��/��M�3�ޚ|��]�����IN5����Ͻ^(8+Apn���ͥ<�4e�d�N�X���3��ϪvH�:��q�'�������w�y���`��pĸ��`E -w������zǞ`=���U�.� ?Q�'���C[=wœ������/3�� ��n���t�7ۑ^�V�?.�6m�"��g��~Wq+�淏Y�$i��/~@2�3VYmN�>ٮO�@����%u5J����B~U���X?��no6x�����S�����rz]�}��w-�𲈦��#��jEc!T0�<Is��K������w��]e����P����&s�Nn�ۣܣE�0!X�ݲ'�?��"�x��R���3v{%YW-k]�gN������/��QZҫ%���3�0�U9�]"ɼ "�&ț�yw�I�%���f��;~-{so�R�n��#ɣ�
��DR]����jY	a�|��� ׏'�+���g��ƛ;�,����`K��`�u>�o�m	; �gCuz��Jr�iem�_�mdJO(�8~���������K�����f���w�o]�ѥ�`�����b�X�_5�Vy��,,��;���һP�����H�(�O���=���P�h�c�<�G��A111{ �8K�kD9�X�e�v��J١�0�J��/�b���y:�L��?~�t/-^��C���>���=��N�h�B���iRz��lteq�xM���w��!��|<����(�!�߽��ؔ�<��{���J�@:?h��x�SR�Q��r��b�l��R��a@vv�ſ��[$BHڢ�>�Y{L_9�i�}��t����N?�R�m��q���*��xz�j���Ug�ʵ�^��6v�\��P���ĭ����!�^�'[da�?c��|i� ]����7�W�S	���X�o�@f@�ۼ�َ���Js:����řw��c���u�Z����f�H��Z��g�G����z\�����G樤�i��8��R��8L �n0&.^�t�rn�(_Y��� ���&�p�t	c�H��aLA�c���h�Ppҿ�Z	>e��1�����^_Gj_K壝��fZW�3K�%/<�֞��H��g��R��SiIr�~s&K���w�}ԭ,����_T�?�������Yg�d�򦺽��`?Z�};�&��2!C��[�|���.v��j2���v
�ƀܿ�c��`;uC����l�E:6��X��EP�yI��<M0=�a�1u�^B�:�
�]�AO�j4~8R�]�R>�ɸ�/Y����[�Uɫ�kj��r�����SH6=)��VXFwy��_Y�p�絭d:���P@h��ܷ4&:R��*W�~|�"��.WM��,�6mmo0��ǬX?-:S����(�͘�����,x�2�n�ݟ֪V��y쳉�*AsX�����I�!�s�sdc�4D��8��u�?��l�cm��w�ɐ�C�=<
��p�:�m���1���J���g6�4�� ۔�߮m��E�bI�~�=����)h��5v��m��c���hp,�v�oH��'>.|Y�,�_�{����<	�_�B�����ݰ��ƴ̯���a�GM�r�������
!`�)y�Y�� #v�X�u׌���J̿�ÿ:(�p�Q���_�M��o�)��i'!����:�����K����\h���{�T&��g5�4_�N*?=������d=�w�hD�ja��h��b����I�+���d�QN���W�M'�m*䘭�^��v����q.�ø��4��=<����]Y�O�y�S���A��$H�0s�t����֒bb�������Y��ec�P)����Ɛ���j�]��'���V����?�%�?���i�_���p"$����!�$0C�3�?H�6��Lm^c߿W;v�������Z�Pwnm�Z�/�,Apgh؄��B4y����rL������ ��j�9�H�g}�pđ�9h�?&���oBt���<|_����å�	��#���1d�[y�I��H����
�N/���n���IS��qi..ZkߚG&����;���H� �$��g�'ƨ��l\��Y-h]?��@�b�^}d�+���j�p܊�V�aD_m���W�>�����2����E'Mq����m�q3}Qӄ��� ���A���te|g�l������Y�>�}a��CI��������!i|q��7����<.$C��:op�_uT����^+�R~`	큎�+W�v'�Ww3�A���֮.�X��׍�(!hy2F���������U��t#�n�9� `���T�j��'�.�5��.�?���֥ n�����-j {���� ��|r#宜���eO�{v��s/����(X7�OJ�d�8�S�Gk�����dd���~T�+vmDk-51!��$^����{��}~�p/�}~ͳ����forMⶅ/};�������)�o͞�����} ���sm.�_P]��C\��?(}�����6V�<!j�1���k-��~�ac�g��mĜ����\��Mo� �\:m�B���,�!�I�} 5�������&u!w���1�p�g�򭻷X(rP�vR�CY	%��_�Û��c��{��=2�������A��1{ַ�7e���,������
A��<�|��V���1���M��+i(�hO����X�߻>���",j�� f��w� C�����Ea���d����cpՔ�54qE?6Xnq�$�V�@�VS�a���>�A��$X�W�g�g�3O���>\��ayr���/l�(�Nl��4]�Ѻm�}�P�l�8�4�c���$��w��,=qJ���u�qHU�~�j�<��씍�9pht^�=�r|��l��SR�I��o|w���E}��]���P�_�H���Ò�g�/V����?$�x����P�_qӫ�3G���wMM�:EM���fe��<&��4W��.��C븠�ӄ�Mo6�J�a/S���UN��Cn,Z�_c �']WvY����]���Z��')a���u���U�nN;�l�'[�D���1>t�1�bq�Ik�[M05�� ������١�ˤpZ��S�O�͐��ԝ&�۞P���x�d�ܝ7<� �[�٧�	�<�&��:��O��&����&�?���meV΢��EN*��t��8��_rlo� �P�M5�`/>���ȟ7!%�֭��&I��O�Zڱ��kv������z��єq�:%c!Xq-C��Ƽ�&��^-����������P[���c�P:)���n���j�3)��i�V�Q����u�Չ���甕�S���/�v���V�-K��/<v�Z)� 
��dv�qR���e��Ƹ��fW#Ww��6���X�\[/D9/����@4���\%%8��| Ɵ�6���0�����<t]�-�����W1UJ�W��hsdJ�θ���鶵҅"B�ܱ�G�a�>�Y� ��I��0ވ�3F�2V�������7"����>�:��� {$!������/�f�9M�$����[�2��/~���p-�Y ��V�<P�e?ٮ.f�\.z�vl�?_�d��X�Dw���5}��-�ݠ@�x�����d!�e52��)�y��U���t#>��./�B�s�wt��a���3F��~��$�S�Vm�v��5���B��ŭ����Qi>c��O�8�!'��A�cނ���v|I�k�c�|��a�t��i��et��D0��O$#�f���`��:Q�Ъ�3i��c�=�<ѻ{kn�t�|B!�V��le�٭��;
�7�]S�C����$PxBK ��������������/������Sss�ȫP=�q������� ,a�r��@Oa/�TA/���b�Z�����{�@	v,N������d�Pˎ�����h��D](hA�6���=�j?qߧq�����_�
�\�*!�$��-��C罼��!�� >���%T�?���1$ [�l�	*�Vr����!U0d͗gV���^(�|q�y�_=��Nt?���6	m�����1U��Ek�^s?�R'WH�\�<O��RQD���>D�J���=N�N�Y���+�'t07��W o�7!mO?�\qP� ���ϟCK��?imA�<�����%�/*�AT�z� �k$Gi }J��� K��4�Ջㅱ-P׆��+���W��ȣH�K8Fқ7>�MbD\���Z\S�R�N~�Q��~��SM(!Wp�M)��dIѾC_-����R��C����;w���� #J�D��v�DQ��q��0��s��������S=����G�1�9.B3��F�O\,..'هC2��ՕI֠zI�sK�L�����뫲ذ3��f�������s�+��)�N�N�]����j��:5������;AN��86F�TL�y�����
h��H��]z]DB)r���_�����Kcq�: ���&[�M�^�c�d�	3��Ղ�)����]&�����!k���=������]��IM�I�a�e��`sn*�Jhm�(�~�N���
�c�������ϞO���}�B�#2�=�N~W�$�*5�� F>莁��<w`;י̶v��� xG����|��O�1aczp��Sp��d�i���p�cj���.0��?�I<t�T���ՑzB��G0Ǫ"�2��R{�����N�F�y1ֿ�
m�n��@��"���o�V?�fص�Yt�e��U�L}�$���3�9c�ȝv�= ��79;ɠnN�� j҇�����	��t\�z�������uA�u(A��
��c�SA�8�����V���j��i��ɏt|ny;����^���%H(�'�\�D��-�����9;:u-���{�������?����'���޿�g���]�3�wj׵�y�2\��?�\T�2M@B�7�!����,U
�v8e ����kB��㶓͜x�?����! t�%zv�,���I�<V+����W.�֕�-$��5�D��+�"�ѐ�|���{�f/S��Ι!P�)� 4䀖l�v~s��t��L��ݽ$��_-
sz��&h�s�v���c�ըL�c�0�G�{0^`*�d|��X4N���\p��1�0$��?5��Ӌ+G�F�&����x�r�,�/��EB�ɓ)���?(@��E��Y䚂��as6�P�P5-ܶn�_O��R�'Tv�����G�z���Iu�'C_�
U*3Tk��k�][t>��uٳ��ʆ��R�]������'�B�_�p��Pd+{FdZ����z?�������7�q��9�
�����5U���=ϦL��~���L�,d�<�,����l\=J$�#��V�^��c|<4����Lfw�:�̎�Z_轧J��u��]�==0�$=�f�����.'��������Vo�<s�kq�b��xM���0����s���� 8� H��6t��{b���ڏ��	��Ꮥ��G�����)w��N�k8��[4�Z��R����#��Q������r�*��Ӡf���SqQ8�a�F�����B����%��X1�ZN�B�x4If����E�a��7�ï��. q0��r �� FHU5�C���ܴƨ�w��7Mx�:�V��'���c����/t ��b�d�_���@=�S�{^�2�;uo�q���/�}�{�hǓ��[E��]�%y8��|�Lr����xuY��Aа�6�n�������'��l/½m��w1��@n�J9����Ku mwC�	�?���t1��eQ�VN��I*����.b��*!���k��^���4��Ch��� ��h�����U|�B�5��P�|��kHݿ�%�0������x�T>���6ǃ[JeVk���T��lj�p96�X�� ץHop^�J\<��/��gti�az�P:��mKs^� ��3?�^�K3�C�P�>��1�����
�'\���?+/���2s����eV^�EnN7sBw�2\��<�Ȉ{�� %�b���|��jݑU�x�`DaH\��6��m��ti=<��I��2 9�h�T�`�q�tr�����������:%���/ɺ�Q��9��2���!�S�ԋ�L1�Q�m��-��f;ي�=ￕiPi^g�f*�p�ـ����s9�R7�w���t!B5���ƜM���?�k�g�we�foČz��9=g��Y�I��#�7:v��&��qa�R�S�=}-��-k�o�R�a��2����T5O�ķ�вp��?C��H�K���?G��gB~�]�KF�p�ͼ� ��~��>	���g�����֦�@*3:?bH�'��`�N�,`X�x�W�"q%+n������H!���y%ӻ���5��)q���� �W-
��EشY!��G�i>֟[�O~��3Z��vu�K�ט
���H�
$�*t�A]
jz�_��	 �ܡx�(��q�B���!b�����7����ӣ�O�W�A~��း�c���1������T赫�h��m�"���l�+Λ���;�"�����Q>��Ę���є�X�̇�Ј��;�,J+x1>f�{7
f�ZT�)ˊ=����D��©���4�6�JT�樟Vt��S��4��K}ּ�{��e���CKU18����޿5�m��`!q�\%[/�!�ףA����k �ꭧR\MO$7���D;���a<e��\.��\�󺶾f�(�9�@Z8 �$�-�v���9�M^�b��淇v�6w�P��l1��D�,�۠-6�H[&��S��F �����f-���q4�nǨ���w_��WhV�߾�DE8�+�B>�`Ź{�^�?w'����Od�;�����N�~^ �'�z�lō*�N
�8)�ވ��7W%��Q)�w���X�n��ݛB��ҡ�����"m����S�}&F�9f�"����d3�'��;������Ƈˬ';`�۬],����G���҇"�I�J��;c������(MV�.���V�Ŕ� '����2g~�h][�(����ܱ�I�P�+�̉J@����_�Lu��J���O���?Jsv�F��r�FS�Cv�6�ەY0Le�E:�Q�Q��1�:/.
�6��?����R?��_��M%�k�Ã�����P�9 ��s������Gt��Fߪ�s$�bp���0��l���7*H��KI�Q���7V�5�GOkL/-
;3�n�h��?���<�9���q��uӸ�P.��-�w�	�xu���{�[>��.�<2*����Cr����P�/��"��"���B�XUa��� *�����"5�̮���ݛQ�-�B�5�?][���x���u�0�&�����̈́�*�"�g��|��x\�*�I�;���!g�>n�c\F�?��M	��:��f���;��Yd��e<���V^� �����I��ל���?&��ڴw9��py�k���a�A�u/�t�3�4��7zw���SgXwD�7�z��ʸI�h�Ј�ـi�Diqr�ij��9����㘩�����U�q���T��w��L
�W�h�v��M1�;�����>l���;�x%�Ɛ�y�vh�aS�S�=�(��(o���g�i����i� ojK�����L��AW�,fJ��3')ƛ:`t���f��s�q��3u�&�aC��O�}�R�U0Cb����)Cuzʏ�f�x;�uYWTQ��ض��u��ϑ ���Z�(�_w�Mf(�P�^��v�S��W�,��	��wӇ���������p�s����b$Z����'f5��V��>�9v�,�1����������呃B�����-E���o����)^�Ć)��9�����{;6@
6�0Tu+4��-�K�l�7��~���Ӻ`L�t*�FR���95x��v�hu���wC��c�E��"��7^8���r�Np�Pߩ�mɣ8��wz�e�����Z��:+Z���Bq��/������-h(�'٨�8���
��U���� w�G|`ӠԿ'|�/[�m���7��lT������g�X7"�r�O��^ ������J���1U{�-���{$d|��8�@ٱ�zu�o���B��g�U�V˷�'W���V9��{9�����T٘:���&;a � ��t�%ߙ���͉ކ�E�l�Y�ҫz�^���]i�3͇�c��-,��/��P�v�Z4e\�p�w維�Zp�ֱ�<r(��~Z���{-����Daﷇ�������Yg���r�ɬ��<���N+>C�Kr��%���?�]���}��J�o�E����&9@�(1��֞j��ͧ�WWl��fLVw����z�N�V5�����W{���i�D~+�?o���Zn�X��K�O�lV��b�~$���d���[��C�A���.�>'ѳ���6�euɺ\�����%�w%��VLK�s��g	��V�s���a��$������~��w�}��n�ii=8}���2C��� ��v�����B*��ǱB�V�X2�� ��{u���x�{��]��V1�������"��	]c�OH���U��������c�t�Pe�;��4�����j)8���N	2�O&מ������'����w�(����l�&��
���}���.\J /�K��x��;%�������r��
�el�&/�p�$� �J�HD���K��V��G����1���y�������[�q��כN��S|aS�*�bS�5���V9FȜ�2$���L�!Ĉ=<�|�{�CA��Z �C2��z�x��b����2/Sʙ�5��/JT%Ͼ�"P]F�ux���a�8���(;��b��yA�Ot��U�����>� �EX/�}���}9C�;��ٍ��;�fR��G��ܵe��r�j��vN����7��m1(��Oap����SJ���	j�++��l�9� ������l�PE۽}gp$���6C$��e�g�����_gQ�|Sϑ�����C�휻k�F��YecG�_������O�>B��ͫ6��<�s��WwO��
g������W�f��U���־+�,M�w��nƮ�y2pqE�Ei�w�߱�*�h�l���7zZ�����w���Y�0���;��:�w�'���)5�{����1E�O�-��L��r-
����sG���-J��M��0�z�c.�xsS���筜�H>��}O��7���a��P�(�j��>�ʸG-=7��[r�X�b�NɆ�������ߠB�Om�z�������}u]��������|���A�����6��>����Py<��u8�*�����˸�Q?�׋3I �u��"��_��<��ʾ��:���r1taW��躝�Lg��0��߿r��8�M!eS�\���O���K������~�կ��YQw���#�@�_��m�'+�!���-��R=�Y&w�d���`��u�]� ���(w�.��ϗ�<cx�<��'gw� ƾ�#�~�\�����҆�;�d/���>�Ue�ʾ��˟��A���,���`i�"��w���R��_6� Z����j�UB��n��d��!��Mk�.j4ew��c)��q04�������?~޷ֶڂ�L�K��p\��%�����#�0i�KZ���e��K]S��k�� ��p�t}xQHJ67�]�N�W��?��IӖ���CQvhl�+��<j����ɡ����Y'�z����\��|����ٞ�Q���)�'���s��#>��WH*�B�LPs��g.�rG$��*��;�'-v���rO|0��Xv8�(����Or �TRE�f(���|#_��~�d�oϖ뒞�Q��� �rb�D�ٺ����Ce�e���˞;�P�T�����f���m�6�\����0Ә^���d.�}\��9��Uk�ʝߡ�]�t��GNK���K��_�M���Z�A�u9�i��M��e�K��ip˘�~��2���B���(�麳-w�`E66FA�J�daU�I�&l����X��|��v�80t����J�ɡJ���]�S]al�����g�d����E:�{�]D�����~�3z'�|Ç��EXfA�_C*������t����6?���	%��6�a��u������Y��#��^#[��<K&�.�d�V����E?1�b����6�A����o� �������\z�L�1U��A-�g6��ح4\�,y��z)����!	�*ť;>A�������9vbpk?��;����|5�E�2�/�z��%��u˟��^�<Ӳ��!*y�v[0��Kgs0k�>�~C��wT�C��V��T�$�/M#�͸��
Oܘp�n4��W�����S�0���P�J���jC�X�n3��^t�M�Yr��+������\���挐�#����e�VJ��,�*j���G�o����?~��P�b��/�V�K�[Ъ:)���fmU5�Rb֢. ��G��N��y/��A��VQ�O(�n�Wa�[RF�g;�@�X�}x���Ϯ���"C��|%\�8&�y'�W��e�|�@�p7dxQ{_c���Z��:P����S4&R:!��z&-�N.KvK�6uY!�,�3�V���:�˴FB�!}+�S
^����Ȕ�s�"	ϻ��{��)����1��K��sSr���%<��سv`��eړAp�=sy'�eQp�oh�(���\����V����t=��׉����K�TTl%N��m#.ÝH~x�f�̯nǭ ��83��UO��Iz���JgTi������N�޾�A;j�L_�O<�3���vump'J���u"��{w�b��~�В�V5�y���[-����g�UO��d}5 �F�2+�R�o������x�4� ��T�K܉��F8��or9��#es��ڬ�4*���'��6���x�Q�z�O��e7�
ӊ�r��1�be���;"	���D;�Oܕg"�F�F�T�����?;6A��QV�f�U��Ti:��>xx{����ۣ��ܨ��i�&i����h.�4l$�0.W��t�b"4^�#�M�@��i����E���|/��pk6it]ul^���A4˹�C>�Bԍ+��t�FS�ohJ�;�l��M�ù���aimMY;y�����5�]�u��B�x�z��S�g��.����Қ����u1���v�^ޗ�����q��l�tlx�*��V�'
��+k��<��;q� �%��:��݉謙�ļZG���F-� �2m�P�i��,�E��/��B�|�%����f���_�߁��uIyO�w#V�-:�͠,�ES�	/��s'��bu\�g�6ž�o�a��m+V��J�FڗǪ����������)DEՍBII�o��a;D��2v�T}���4�b��]�O�n���-���]9]�V�]&7��^?2"4�:	�ӈ���X�i����,������cU\��MXUl-xh���=_w�y��Ŏ����Ӛ�孾w"����͎�嫽L�Ew<R��̦��v���������+��C{�z�k���1���*�k=]u<��-�3���䥨X���a󏕜fSy�3O!C�s������Z���3dK��8�*�JL�^��b
:z"����[x����e�|��6vׁ�h"�=xF}u�=/�JY� �w��htVLkT1s�笇/�$�����E7�,�ZqpeE^���Xu�=L'��������o��Y�<�.�iFH�j��2 �ۦ�4[Os�ԓ��Ӽ��P���)Z�J�t����㟑TŴ��-*���3� mri��/t��I���p߸�������XY^��zѶ��T]=��oe�UT��y3��]�'["�%:r�����+�l��#A��NИQ;�l���m����>�����3HMn�璣$�{�c���OY�R�Z,�s\r�Uvgmj����� �P93;�7ɝXK䂪��*�a�L��?+���4A��W��p�g��Fx�ҳ�z)ttu\��g����d��U��Kہ�H�i ���&�]S(ڗ�E\s�JWj�P�'��=ϕ�X�6v��
ވDc�#wm5�����BP��xNI鬌(�����gn�E&�Q��=�l@5�
=}*6IWm~���3 �Q�T�8����y�nŪ�>�Lzڬq��M4��ɍL0J��&s�� ���[����ع��.~T��[)\�P����jM��`'X�G]�'�#�iQ�*�"��xR�úC�'��F\=�:J�O�D�=tG0��ܽ�菧�n����DÒB��5Nh�5�e"R���K���@~�yKR��V7������d��V2�e2��|bF�Z�f1=\�&S�x3ud��R����=�� �Rْ�"W�Z�^Ox 4pi�+�3��*8Up��'����X�ƃ�vl�r�K��bX��_������<w��^'^Oό���j��>��c�&a���a�IŚ�|�]�z/�{ȃ��7%�K��́pU�A,5	f��O}1���މ�X�˱���}l�<���W���J�����
S�N�F"t,�Ȗ,�ӱ��0�X��pU�K����+1���A��Hgl*�@��{�Э 0Ah<�"��,���x��7�޾sؼk�O�+��;���]�uu��3rSӰvY]��/�ro4�0��XO?�M�Q�nJ� (�x'et��� >��G�[O�[�]c|���0̀ܢ&�ѯZ�>w�%Z$��w� �Y!�	���2f�I�V��[N�,�d��+V=1v�n��)��u_t'�>O�p�g_�w��M�Q�^H����#��.�-����iI�����x�b4���pyVDC�����aMYi-[������:g{"Uq��ee�����<zO��ʪht���)n�	T��͞)cV�r9��WQeη��T쥡[i�E�wi�SƼj�ba҃3)�����+�hPF�ɖ��|f�u�~UO�j%.��;K�FM�"�çI&� 4��F�j8n�P�w����&gw)I�N���j"Yq������.c�*1�_&��*G&nx���˿:E>�z�B@_'>��]J����f�k�s<��w��H��:�	ַ'b��>W�$]�j�l7�&��aצ�h��<��׊��X�(��v����6P����S��Q�eNώ�Ό��;-�v&�1,?���y��*�M�:z�m 0 ^+U�ƽ����:��$@�,���f,�.a�;�Z
��y����%�J��T�#{�x�mQ[��K�E�ci_�n�S!XKjϵ���:ǅT��Up��_��<��h ��x��ت�J6~oN" �xs9�AK�:~�^���e�υ���4KV�����V�l����1�'@����R?�~gͼR�xPO"?��K�e>�n��1f.S/���,�J��Ku�jEUx�����+�f�S��<R�'}4���)L�-��;&�i�h$�
x)���>��É�a�@���w��7�@�3���OA`��q�xI�c���Jo�6�2�wЋ��s�@"E�����S����U0a8T�sJ*��~h�&�b0r�z��-qr���t��?!�pL�ͺ�!��'��N��qka=��zC֦�c��k��pƟ�#S?Tߎ�A��-9�[��U�Ö5�.*��[)]O��M ��8�o���2s�׎�-��-���~���燰[��C'�U?U{t����-u��ݓ\���5�S	7au��"Ȟ�k`G�{�V<<-�٘���#��f� A�!�c����kz���{"|~l�Q!wPF��H+
���P:E��>�K|����>&v�ʒcۭ�>VJ��ߵZݙ[���U�|V	�����P(v�p��8�n�փ�YE�퍕�؜Tԍ{�D�	����V�������݉ �LI~��4���Uk�k�{.�NJT��qY<��<4��Ѐ�bG�*�		�2���V�k*�d��=~H�*z���H}���@,�� L:�}-�^8Rz�r�w����*��*=�/+T�h�5i ݝ�e�䪙w�����R���!������O��P�5���	����y45��/�8�b@�z�` �Y�N�2bƶ�D�b�Y�a|I�##z�����b\ª�v���4��4pĝإX�n6�Ղ���]r�Y���z�*�4�؋.�b���_��t��
�$��{�O$	��+3-aV΂g����9��.�mi��sl�jP`��e}�,I�~���W�h�Z��;�8�g��?�����@5���Ý�����Ǭb쿉n8>���ׇ��UT��<��ii>������w*�$���Kaq�W(�(���Hگ�/�J�)�����[�/5k�\�x|��$Hg�RT����D����f;A�e�K�< J���� ����iX��B����\Y��� ߔ���hGr�t�4ZP�y*3�i��c��>����ɇ�V�4�1չRp[�A#P�`��H�T���%��VD��>Hݏ������{˗���^@O��[-���G�q��$(�W�.t4�z��DJ`?L�!�j��8@��*�XżE]gYd>���e���f3��:�#O�k{_�7���p:�:2հE{��j�M�Δ����/�v��C�0��ߠu�~���1������Ӥ��+�T��N��ҙʢ;QO1= &�5(�E���5u'�/\�.Rm~�rW��C8+2�Y��o�
�.��[���Qug�:9Ax���F�����BN2�i�v���r,ҷ�fD٦�
	ئ�%�a��s��L&\�����6�FVS��zb�F�	�/�p9\�0M������G��m���K��bƀpVǀ���;H
�nk��^8;�bW�X�V C!����+O��l��wp�n_Qc����ה�m�xT�$�����O�Zu����eG�>�ܽNa��.�wkٶG�k"�='�R�s���	L>-)��1���&��O��"������y�PS��r�k��d��gbC�2�h�:.��h��w�W�����۩���;e*�V�i)�2@2�wJS1c�r4c�>�qv�<�q�c"C��L7�j|X��S_M�@�lmעo�����ċ��f|0���Z]}y$�_�΋��b�.^:Y~��?Hv��VɈ�
�fh|�� fxe�p7y(={\̴7���JP�J?4���x&4B܉>�W���-H��.���]��sKM�T�.,=H e�jd�
/;H�f\�4���*V= �r>g���n=���Q!�+��e�jk.��1��,�4�6�Bm���#� M�)��������F���?W�RN}��c��a��k%5�"yx <����H�*$�bǈ�*7�#���wl���Չ7`�?�WA�����-��q-u4�4O�$ϯ�ۋY�Ҵo��Yj�^�0��"��m�GCZ ��}�u�cOAn�["j�?Y������Y�U�(R�+tѕ)MC罽cz� �g�.�*w�3�҉t��5� SM9~�p�ݔ3�X�)2,�F����S+�~��\��,`q�	B!^����H[ K�i��_��EB|'9�k����C�Ñ`�N-y�ꥊ�ȻVV�nQ.�,�0K�W�q/"�EX��g%����.��BM��s6�c�s�͔c��O�ҙ�:�}>� �A͔�M�9�t1��̭}G�҆\�1��d��%�S���D�x/��+�����h.�
�Y|�ұ���W�\_�TM�$�؉��A��dk���qG̞u�dh�u��#-��X5�R�ޥ�ѩˮZ�B�ϊ�yY�ȁ�}��e���?pY����Do��#�Fd�����)fG�}�|���ɬ]D�X*6��d�{-(��x�a ��Xj���ైba�
� ��2���͞0x�ԡxڷXGE�,; \YO`΢	�.�k���U�;q�&1:.oh&���WT��/�~}q�����.1+�]
oi�\:�e�8�4�Wi?�*�%�I�陈��*�y,�tZ�σ/�g'��H4�p+���!7^��,r�R���"d��m��'6h�$�t<y���W����a�����QG�8-�N T��\1 9G��K߲_���g�����zk����yj�8E x����'y"c�}^��#2�w.MJ��c��J9�%�FN�JX�'���\$��:I0Z�)��0�azg4Z����Х6|��W�	�W�L��!���
S7�k�*���:$̝�Y_Xrh\_o�]��e��d����BH�� �8�!��_�@��1먕�l��NT���֑�rm��&�DM6��ęj��eI��\m����4r�Y\�NpS�(�]������a>*0����8_����������J�%Yw�?t���'f㦖���9
��>���R�B�iP�J��Q�.@;��M��ef��r�lE��b�$��n�(o�QI�ud��Չ��.	3\�kc�5�rƺ�a�`�p��@�=bt鍁�������~O����un�31ݛwY=�@7P;XN�v��9 ���w�������k��xO��{�>ˊ�d���X��P.��Wm��%wө��'��P���
�Bņ�2�9A�4n�=e�z�>ۆ���rͨ�B�:
�V��dYx7���׹�I=���Qa�ΨO_�!�z��j�D*��R�a�����p �zH!����,�_���y7�C���'�N�&���q�>g[�"��"���W;�hۛd \S����2�4>���q����u�5Tu�$����q��F�jk ����7����,�j'ϕ|�{D�n�7���k��T����^���I��YW�9#���E�PR[k+g*֮�Soyi��3A0\�]G�N��)т�HBݪ�1�
�;(�u*�bK��&�Ca�:��Ƃ\@[͌��N_��RZ�(Zp'�&�4Ԇ��|��5=��,����C�I��z̀X�q��?�����
��Z��<r��1�����ڳ��N� e�WT-Z�zωy�b�s��+|�I�U����*�qV\���|U�"��f�+�]FmRd0��%��zJ��y�7�잝���;9�W��sC�(/D� ��ɡ8V�`J����*�_�?��wi��[����ڳ���0q,�����"�'�k���X�K�H��_R�>v���!g�s.iJ�`b/!�vf���R�����X cZ�U�b�&Y<\k��⦭�_V��.\�0p��y[l�<�k��މ�͸\vu�||B�*s~~�������Mlnl�U 7�Y��/�ydH�٧�<�l�$�>|��[� ���F���Dey?�?��ӉW���UNgq{v���Z��茇ȂS]��H����RyY�o��~	�T�`(SCW��yo�.'�t4��j/�
��,�X�s��DU�f<�]��'�0Iݸ�}:���'�n��)[	�%�tU�m���Đ���޵F5uea[�:�mg��Y�ʹ�PS�-���(
(>	�X�P���bY��*��P�
i
i*܋�$�y��r�P^1@��!�I�KmWk�8�5?{�%97��s�������9 ���i�m~�P����}���D"������α.{��03���&5���;��7�WuZ�����N߹�!����|i�����*���R�]��C���i�5~��7�9����x΀��t<>	�t ����+^_��*�8��V�W_�߾�?Z�K�UG?�nP��_� ;Gy�ybw^ĩXֆ�\0/uAW��D|����F��\#pEKֻ�n ċ���t$kq�(���Y��5C��d�֏D�?�ֵWe��� �yH�ATսQN��%�x�}��1����a����U�Z&��]������[7-�~�SX�����e��`����}���5K�g�j�g?9¤m�?�|�C�ǽd����spNy0�;5�s��K7
@d�~N.�1�b<��V���d�Hx�/������B�j�����uo�f-�Mӵ	ߓ��,Z���v�{�rg��Z�^t��7��f�]N]�<�1c�Y>kE��`:/=9x�ż��܉��[�c�s��ַ�(�P+r��.����Vc�7�wvb�=���K3W5�@R�.�"%?����%�=���MԏPzw�TL��B�U R���Uy *L�ߞ3;��w*V��ȍ���+�7�]z�U�n�������Yu�fcJ�ԛ�@��o��y뚦` �iE+[�窮�l�q�4���S��J����LN $Fx���"�c���wk�����y��z*��hZRJ�X�G4/V��L�_�X��n0�X9��s����A�V?���@���XEϱg��h�����~sm�7i���S5=�SD4�	+6_�i�'�&�!�}#��K�g���W�]���u��7��5Q�An��c��!va\�H(�� ҄��C:'�F���OGP�] 0>�H���l��)�i!���pz۲�qb�����CW���Ǣ���9 ���ڊ�{ϭ��Z|���~���e�q���@���\��veO�e��N翳��`4��7O����rZ��9j��*>�m�0�f�UwV��ŵRYo��1�ڲR�Wy'~[H
�\��4e`�Ё�)�צ��M
aA2f�Y3EqQۥ�<Ǐ:�1����M�e+�y^�$��=�Ĕ��}�Al��p����u�Jm�4V��?�n4JF˽:�����d�*3�Q^�40�Y(��m�\G�ٻ<[��޻�s{eX��=�L�s��c��3~w��G�ǲ�����c]F��WjIy�fې91⌶Vy��{H�1)����uPȰ�K����:ld̇��IF���O��0����|�h�փ�r���˴@D�e�6��e����]|Vu��\U�%����:��7�y��~�"��n���Oǲ��1k��#%/�頝!��El��lZ3a3�+�s��I"�28ܭ�?� �m�	X����T=yy��D�#�%3�m��@4ec�	"���P��W��� ���aQoH��(Mt��4��V�i�M2�Z;�PG�ڇ�a��2k�priD�!
���=��[�jq�	���!k��U�D},��Oאt�P�%RpB�h����c���s�H@����7���z����H�F��7��nZ��HdKO`��u��O@��]�YLQ��)D�U+��BMX�����ION�H�S���=0�EX1^l���5���m�FW�u@��[5�D�Y1%�U��N8%\��;)���a)g�PiG��s<q�V1��kG!�,W`�ǲy�2Q�
6Hd�̍`�Z`&1�p�{���#�̡ݠO��䶾�Uȶ6k�n�E�M�nI�$��.;|(�٪F+�_�p\�Hӳ�w���祉ʓ�F���U��NP����r&����z��#n�#��d-�,%>1ŧ�3�l{�lOuCYbe��^I���L���b��T��'$K���r�l��m{<9m]t�9W�ɯ�g��CP{��4IZE��gĐ�u�YD���*x�3_㔬�6	3!l����bvy\�'�Xx�t�[���oZ,M<�I��̈́aC!�z���7%q?(䊾:Eլ���C�N�[Z��5��C�����f��CQe��a�b�N�����	�(���ڈ�U���v�m|��A[�:LW�ȼ�zQ&�3��y�7)����TX�x&Z^xeG��Q
��]c`X'� u�tJy�-F.n��a�����-g��o��<H폔	�T����e�_��.)g56H/8
�A���ɼ��,��ٱW��n���{��$a5Lr�{�9�Q4p�l,�9���F"!�<I5����-C1�T'墪��ot#n #n{xr�v�@`'���:T��A@��e����U��"���Vv���q;
3,K�&:��E��w-غ�WF�5�8�Vi� ]���n��݃g�]�
bP�
3q0�gu�=�Y�"Q&�7�����a2���ZB� �0���0}	m��{���m����S�y�欁k�g��W�ݛ�oPK   ���X���<  -  /   images/988d5287-ee6b-46f4-9561-988eb80bd729.png�yeP^�6�t������?Xri�n�KAXr���	]@b�%�N�K��$EI)A���y?���;s�s�������M6�פ"g#��ã��R3�G<<|~R��}���=��hY���q����t75��d��[�L�_��\�Eݽ<��}\E��^"����ػ�� �A���i@����-Vl����W/��W�+L���j�(�o;�?\w��2j~��/����6��ͫ��&�c��(}-UJkL�؋�Q�r���K��_M��U������'�j��u�Je�q8���|d=N���O�E�^U���J~�����N��륞Ў�0p�JmKK��z���B�f�n1���c2|V�B�Ȼ!���fX�	����p�i����L�QU{m�a���,�����lvv�Ք,��@<�*�#��/��зYQ�j'��a0X��mY����~MdJ�C 7��%CB^Vz
�&�)=�����t�%�`l��K"
5�n����pkt$E�������t�N�eO��lV�&�hr�x>T�j~�!�9L�TN'yf���粔M�M��M*_3O�I�xU�+-c`��\�dtdd��D�#u�c�����҇ۧ;�N�!!!�.0XW!�8/_s7?oD �����l�N�b���V��2�ŋJ�`��	v�=m�>�Q������r�-r�S��5��o�~�:
df���;�����������J�~���̓�����r3U�[��8�DҀ׺P(�u����Q��[�������N~�v������(��L���=}�CAE�r�P��tR�}ȏ�/�b������v<�]���6�Ă�#�C�1J��f�+�r#\�RR���;29���/�������t����&���R�m��_S"�,iu\�e6��&+�ᝉ�b72����J����3k�����:/�'���?�	�����ީ}ĝ������v��'�);K�T�ͤU%��"3U���i�RSX~'�;6g�%�Y����ȫ�/��{iI�U|�
/��rn�P��랭"�Z�=0���Tǫ<L���qp�����R��A�Qd�����q��렽���/\MUΞ��"�ሌ�5��4Q��U�ھ�2��}5�J{�E(�m�����=���4}m�����CCC/���rX����˝�U|�D#��=�r�,,:�~���y�6*���gnV-s��Y������zEWb+;����Z���`E-Hĵ,���Q��p��V�}W�{�J7��b�e�B��'�q��6�o3,�L���ә,�ZBP*?]�uF�e��%^�<ӷ�����0�w�p%}R閞$ڿl#�^��k0��V�Ϝ��Y�����<n�~��%�L7��֛Dcs0������>\����ܛ�o{l�uejs�Zl�,�?7��3-=�;��6+n��T�bp�]l7�6���*�q[���0���'�\��ͅ�r�3���K��)������clH��Q�4:�,B�ǂA�uO�:I��&ӓ�Hn�s��fż��5���鴀�����E��WwF/�jo��t?]�j��!7r���.O ��a=(�W �k���i=m+�"Z�7SY���l���EJ~$T�v`���p^7��{H��}M�����f�� 
 0�i!�h����u�|�6����e�a�-	U���5�w�NľN�Y@
K��s\=d��9�B��~j�:�t4pdz�MJVi-M��Q��y0˪��`�⪣ߚ<疜���?�y�I�RHHF�ODd��;&<炈R���>e̝�����x�L��}c��0�4�.�gY9�z�h,`ѫzT�������J�3u�/Uf�����������3��ExJ��o��*�S�I�%�0sw�=���<�%H��G�l��f`	�IʏKK����7�U�qw�hϚLؤ��s���>���Mf�bƎ�-ﺍlW�NX�Ť/[�᫫N�~�0��v��3
�_��7o�K)�3ˢ��N�K��tw�/�{��:"Sumј6"��zC�:�@Wua��?�}�������()�L��{D͡d9U���,2�O>����D�Ld0��Aϐ*744�f���FJ}��[��)��Q6?�����-�|{G�w�\���t^o��eM�u��#T�Ҽ������a5{����Xn�wEsƊnr�̒�-�pZ��~�g�I���G���T{0�~������̒L��H�����"ګ������O�����GMk[��������f�%1��Js.\��s{ba�c[IT��
��`�j���s��rz�'+�'EW��5��!N�8�� r���T ��C���ؚK�����z��3`�[����W���@�bt�;��9��~(�Km�`afț�D��
zM��SV�)^��44������Qv��2{bk����y��&��|��.rj��t��˻�����g6z��^��)���	����~��tM�tnFV�p�,����m��ĳ��ج����h1Yp������݂�,���[(��Ѳj�3��+�r�}0�� ��BS7Y+%�� G�j(T^�׃�XM�{vo�w�~\�Iz1��
�l��'��O�
��)��O��8^��za���=tZ����4�@w&�J���\�f�2F�h-�X�GJh���e��&�V���~�;�c�o�Ɏ�N�4�/x��lQ��I��UkY��{����>�a������DG�s]T�=�6`�e��-��kj�2V8��A5%Ο�*�x��a'˚����܆
�|�udBE˒��f�(jOL��*�B���K^�k��?@�%�RBn�<�1���#���fi������T���4�583bCұb��6%���Ds�v�k��'l�CY��u� �3
)�ٸ$��6U2�ˤ�ͣ�b�#v��ѡM
�K�|��^Ir��U%.iЎA���!�h		��ۀ�����{��z1���K�ݮM�Z�|%����'���}~�Ѷ������Tb���z �
˙�={�)AQ��~?�k�j��E��[��s��?a�W�m~� DR�mv��<���@@YN���g����k�T�H�>f�]��e�IA���&��"�J�{�2�Q:�>��T��\�y��GԂ��^��ADg�]Lܬ���Az{%�4�Q�ǚ��(B��9���Z�f�鮏��R�~�Z�@��	���T�G(|�U9ωz�=�6=J��V�X�����{�;1tOI��Y��R�	��47��$�+M�P�YHQ�Y2P�m��8�Z|h�[�T�&���Ziug���j������6x�[p���G6�� E���SQ|��u2�׭A��$�y"�l;o��e��LbQ[��*�ss'[��(�*�Q_��X/f�
d�xq����]g��u�~��ٴ*\.��@��:U��\���Xn����Z�hxp�h<w���)]{���;
\1"Ix~񶠨�~��Mfm:�t:ja�u�:n��Ɔ����	k�&�JQ�<AU�d�����:����J8*������Z�5����C�GD���q��vlĆ����o�\���Xvz�C��t�rN��g�J�.8�������У����T���Sm��nI����z�'���7��K�` Z�����qk�Sߏw�PQ5��Z��&��!k����'��{w{�虑�Qn����g�i�4��|y�v�. W���k����Qݪ5�I||��2e�_�yɏ��~����H	d�aB�=Y����4����s{���Z:OF���8G�����|Q����퓵��c��ȥv���O��x�d'��3hw֖dh��gqF�
?:�����UeTU pq�$��hJ�V1���&�L#���]A�Q�Tb�r���6T��6���-2�U��I�
�9����g�^��\`��dM�~cW���=I�?6�S�4�����ނ�>�Մ�}�o�K~>�
|V�-�E�Ѕ{���T���b�ϰ��{F�8�1��t������ 9ǧ�f���\u9�	��6��=��&\�򀂏z.q����s[�ŵ�S+�^�������"�@2�1C�gL������nv�k�pB>v�@�+%~6%�Q��50X�@ѭI���������l_\wv��Ǐ�~<���n5^(��Y@\Y@3)[�q?y�:<���{Z �.�%5��%%��b��P�%� Ы*A��b�N��]��]��ma1�
g5qj"�<�52���ZZ���a�Q��OM�$�~թ, � �$�@'#u��G��:�[��ġ�'��ԩ�(dL/�)3)�SŨ�#�5�ח5�P�����e{6�L�8��a4iY��)����u��h�e�f;���Ie.����#�U�ɢMP�(�t�TՖ�� !�RR�+���21A��B�FR��_���D�;F0W��ԡ1p(�#����݃�K��-�[�~���TSa�t�0��O�d�r��'B��lid�a�C|��]���F�تa��^���v{8�	�ֽ'���&9��� ͢?/2a[L�8���KB�`�V��胔J	�݂K��� kA�H��� n
ɒws!8�X�����k��s��lax[�U�ϳwK-�Q���v��7
����z㛭_���������N�?/�Yi	T�J2q�C���<|��*�@��=��'�.�=a�lO�����s&Yn�8[<+S�*C琡��H#��]a���h�G���1B`q^���F�T�v�U�꟫�Yd	L9����f�w��V��N�s͑*��tz�ƣ��p�!}����L�s��ܽ��m�Sܹ�>���y�8-W��g{{E�bԉ&L��2�鐌���ExOV�2+���ƍ!Ø:���G0ә��j/:=���Z�D���p�6�rl�wc���K��lZvO�A�����U�W�lRY4�&M�w:�޻48i�R��nzX�����n�a�>:$F'�G�%Z'�d>l��f��� �ag�MG�ߪC	T���G�`�X�'w^�v�������x���ąs�ю�W
/��ٜ4(����\'���U6���S�<��
A�A��z�i����O��=�3�8<���ճH�N$�Y�©��wѤ?���`r�)l�����a�Es�1�ڔ{��r�#3.&\����~��V]iw^�o�`��us�X�Ʊ��޹3RK�_
�7�V��YW��1P�.���lT4�1��Wu���4�p��`��&��j���7:�&��+�����W���;~ t�:m�3�PZl��kW%�X��}�N�Հ�+~�'%�V����F5ҡ+@|l�aO#��Iђ ��,?�랟�k�}/����px��C�ƍ���su�r���aiv�|�B�i��m�z0>|u�ې�D���>6` �A��߸���p?]'�����@<b���j���wZ$�f��X;�brӴb�=&L��l��Tm�$�� ��h�1�k���/h�`A��g�c�W%`����I�ja��)�S��/���Ҩu���]Tep(�^	]�ROR�#K���ޠ  ��&��L��Z�3�:���[������L�S��	:��_�����nT�g�-���s'9ѯ$[bf�"��E��rT��7 �!����p�:���c1�xA�'⏓�p&��0|Y���شjcۥ]���˩5�\�S3��I�F�N�F��#��7�v冬B]�}꛲�t
����kV5�3��GPg�$�Ǝ��ڻ�2����B)Y���'�ϱ��?9+w�{��nX�Z��Rv��쭷V��B��XT��%]p@�E���LW1K��}[�1�t������3|
�1ʰ�P�+�W�d*jJ����a���_6�Rش��g��4�%w���捡v��XO>o�	�!g(4�_�u{z�bG	�� O�'��/�΢I�{���8>���O�M�*] �M���W�R�&���?�#�<�j����=�7i�l���0p��8���>����᱕!�?���85���W|��O���l�z�?K���h��.+��G�ԏjJ(2$�'��	ݱ��J�e�'��a	.�Apg��8�l���P� �D�4]��fR+m���;��}��
�õ��y�!�{�K� Q1;�gO�ɱk-c=���W�O�rc�Y�	�4d����3�8+DZ!���^���b &�����n&�i5D��x�K/�W�Idv��+�:��*�
���k�H<�@.hgW�V�4}�V�mO��.�:�U&��,+$ѷ*ޏ���4�ڋ}e+ݎ�S��^�������(�:��g�����ԋ��V ���/}��7��h�HY����Q챺���E29�&'����?��ـ[Hɗ��f���B�A��$ɢ�d)��ʊ�^�q#���%A^�
M�!cU�=��>��%��n�`��[w���ii~n���b�@'.�>QSB����+b��*�E�A��.�֋��<@�
������9x�D������Ǥ��ŵIv���?���̒�]��8�x����<E���P���{�(?Pou����uq�y��\eE?I�
������l^��e�F���*�jA*�?�����7�sO�O�i�^�G�������&��9�_a0�����:���I����ȁQ����)M��.D7�������zQ���W�K�E��۹v�._��\,{��P�#�S��~ �Ug��kAm:ĳ#8c�喓I���{tIJ��l���@���p?,����s6kЗ|��'gǳi�{`j�Ό�;���w�L�|l^��.K�~�I�4C��cq��M#�ҥ�~��>W�?��>��UIL���vb�R��~��#4�U�}�D�~i�뫡Ub�PK   9l�X�� �  �  /   images/a80855a5-8bca-4bf2-b044-5bb17264cccb.png�l�PNG

   IHDR   c   Z   �N��   sRGB ���   gAMA  ���a   	pHYs  �  ��o�d  (IDATx^��Y�^յ �]�]e�l��`�'�����f0�&$��Cw�H��M�Z�_����_�ɕ��\)t���:�QF�!@@p�$��l����\S�o�ZU��ܨ�w9���k����k��9�2303p|C�X�����O/y��g���ݻ?9444���5����yסC��;:�e�|xx�stt�k��ٮ�����#�ǲ��(�|P
ZC�|0`(�����םq݉��dA�cdd�kV@�ώ��#R�J�3�#q=4��h[���G�D]�?yg'��<:J��ޕV���H�'o+��(�F�̙3400��D����?��7�>�����θ�;��������w�=3]���[�p��
�܇�K0-���b�ZY��GC^��^{�����F�<��*m��hř���褽:<�7ٕ�~��ɟ �U�,C;��sL�i�ڵ7�p���"����7����o��	����ÇKDB%���8x�`5޼y�ʁ���L=�a�y覱�|%�8%�\O��'����~�ܹU��ɓ�N�\����k�<Y3�������o�n��8��W^���xW?W0<F0ξ}�j� &�1dHBe�I�"�'�t�vi�=�y�"p����/��5y�ΠA�}�h�g2@+�Fr�|S��g��l7�?|�W~}���oV��#���/���v��w���Rh�Y��`@ �.G(����B�l��o�?��e���孷�*��^�2�?�և�<���=z��ь�*^������-ep ^�,upB�{��=������0�3|��}�w~����t)��;�Bt���z�Ν�g���£�E�ʩ��Z>��O�e˖��g�`�A
MqB��T~��ꈄTԐ�nݺr饗�ŋ����b2@[o��F��6yɦ���+W���j#�M�_{�cǎ\���領��)��2�w�y��n�d7��B������wh�s��w��P mD4#C�h��ԟ��'��_k����K�믿�,_��2��Xo��vy���֭[�BiNH�@��>��r���|�3��d@�J�<����.��9�g�}v���O|�3
��}��W�� �4�O�6�U�VU=�e+�	
y�u�UW]�~ӦM��a꥗^Z��_���C�1���D0F��?�i���~W�T�cD+J8C� FC����{�n�����O��"���6�F9��j�Ƿ�$?u?���J�U��Sߚk�tE��%H����?���SO=U.	�[�={�Ԟs�i����r:��^��� ҳ��r�����̿������!U�A���/�#@2M�Ҙ���o����p(���HC/�0N3��wB^
�����J�bY���Ix�s�=u���f�Sҡ�����*�\hkw�]w��� y���UZ�5b��4����[��織e0�[
#��o[^x�ژP�Q�9��*
�x��:����-Ҽ��#��ޔ�
$�K���-[��Hf tS���U��ɞ	d�E�{��2?���Z�,�gϏ%�8��@;I/��{ｷ����tE���W�6��3�K*	�ؒY�%�5��F�U�30T��t��p�h�Ӊ �O�`��ի��K��̆�^@ʝtZA~�^�n,�+-��_`ȳ��� zɗ#�Ð�&z�g�E����X��K�E�"��R��	G+��,'�{�h�TX9@?����p�@:8��}�b�t����4D�di����lrnA;�U����S�O�8i���~��1&K5T�e�]�^L.;1���	A�,���A�ɏ.Ϝ�x�־������g���=:dԆ�p�+w�8��>i'��:e9%����g�� ������@��,�<g��ؕ�Si�������|��6��H��C^&��l�%�	�>i����V|x �92!�G��4�\�)��� .��H�9��b&�@�U�@�W�̬t�Hlk��T�QSpEU4�d$��y���Q�<]�ٮ�A@{8 �{8dq���:׭�	dh�E�x�S.��z�9�Қ�'[:\{� �fO�
jE�ΰ�i L!i`�̞�B�J]d���AW��1'��A
�H|��0�(��G�p���/�֨l�(K�Y��'����a���8�)v�NҦ[�S��]C�'���� y�����ke�w���:�}
�z�����G��+=묳j=@'��99'd�e"9���i\�Z�:8�0H�@��_2%�q�峟��x0j���5�\S�����蛶j��O}�t���6
-p�3���
|�s�+K�,����)��@as^xa�(h �_���HG'~v,���Gx)���Z�:�0u�\�{�%R�K.�d|��g:�|v�xsT���L2$��2r_y�夓N����0�hy�k�p�uX�#(��<�OA�����#��!������<�BRX<n�8V�#�KZI_��/}�K�N�m���?{����5k�T���գia��/~��~�鵭�tTʁN�I��Qd�#�>
�ց|] ��a*%%a���k�֝�1/�@A
0�7���r�g��Bk'ǋpNM :>���/ۑ%E1����}��	9'���2��<�h�`�4j� BWO����K,�~ �<�H�%�p�C���d6,9���RV�I+ܽ����tƵG;#��Qf,%�����(d8��W�Z'V��,����z�D�9�S�������ot���k��Gt��*[*�e�s��0^�sr�.����򕯔������4	��&�/����t�6h
\���+*]=M�R�C�s�tHgT+}�{��߻w���bF1BQ���ԍ5�)#���x���Kcen�P?�N�8p���
���r�iD�R^<��*	���.�uӗFF�lIntї���Nr/0��UT�%O�ze��ͫ>r��0���cFPu"[9G�F��VA�iX�i�j(kn l:B����!�ϼ�:��7���J�)�&��<�38�#�:�j/��4ԫ�V���&ߣ�#�����T2�.��epZ��J�S9� #}��M�ʠ�>q�P'���(�w�zq���8G��?�Gc���S�b�=�;:B�@j�R�4��J'@.%�%�����Lrr��à�F�#��1���H�+���t����j�K��1D�i: ���|��_�B[g�I��Z�8�ꌘX>���_L��	<���� ��j��G: ����q@[{��t����s�r͝���#d)w�C�vύX����{u����;ľ�����%/�F��oR�i��v���� >=��=cʁP��'��Gv��8�޵�ܱ3f]�1;�̝�H�GK;�z<�'-��I����j7�6gpH�)�@����k�g�"���+1>c9@����9�6��h�gP����+���מ���<��LN�s��w����,�����K�2����(��x�{�������bwJ�x�[���H2l/�v�m��?�y��[ʽ����=����6{��T�~r�?���a����� �Z#,�A�3�g G��莧9@/aeH�cHx�8@9�
��.��|��w�{��3|o��GO=�v�p��w�?����Ϟ1�Π�������!�8y�NO�v��=�����y��7�5�-?��c��k(��(���R��8��{���Z�G>V� 
���XC�zF�� 1<cZ�' ��c|x"�7>�`}.��_���p́"YĿ���Z@M���o~�j|��k�m�;|�,'�xb}�R�z�������겨�xx,�:#��T�H1��4�f))uƲӰ��|�5�����������T�K6\\vn��������+ʒ�W�\�z�����/��������|}&�9^��x��}Z @<B�OW�Hh[ϰV����dg]�xV0<<Xw�'����9wmMg�uv���=�{�͡X����a֬��4��b��Ǟa钓»Ce��m������g�U��W���ϖU�V��/-;�6��ѡ�2gv����:����H�l�gN,b�(�1<l�;�NI���k����MG��KZe��0N��=tp�F�`,+O=u��|�#���'�<�����t�0�v͹�G+�������6)�����_0>A�@�����-$���])���{�XCۆ)$)�g���cJ���fNVN+V�������������/:�X����)���O��}bV^��0�{�h`NȹFbh�����ϼY�3���ڦ��g@L~�)����7a�8�cđ�� �1u9浪�!c��Y1'�S��H5���Ç��s��f'�u�������\=�gi�]��3ꇇ�KW�<<;���ѧ~���od�y!�<�+=�a�!���^#�����|猶��������f���"T�u4�G��y/iϘ林_~���xQ�?on5��|`�P9���0<����mG���X���(���i\��yu��Q2<ؔ�νg���m��'VS�j)W*CC�˭I�{Vsf�x�E/G�@��m�|n]ٴ��k��}T�z�F��(����G;�|��@=��[�c�[;'p�c:Q����J����|���HgF�?a�ĉl��`���f��C���#=<%�/�GoLY�5��7N�6h���[�v, �j�3D'��O{I�
C2���P��Ә����_9�9�Y�~�5�2ڜ�F�7�0x7���󸦮�e��c�`#�Hf:�}=��ƀ�=��Q���N �6,�?n$�;�b���Y$�D4�?<PWm��a\9���9ti�Z�>���p�إK���vS��9e9d�F��1�m��R?nWo�`���^n���j,FQ�`��̍}D�/�yh��C1g���b�184Pۡ�]��t9@��/�\²�vrm����t@�zp/[ͤ����~(�<)WO^����1�Pa�צ=�3�9��WoГzz�o)�(�Y�'��y�_9�����En�1����My��y(
����+�>r�7�y��>8���[b�|�]w�����{�}�=�����c�����;�<POa?xooժ��9 t���]�7��W����~ NB�G��zku���t@�z���1�u~��m�|�r���K<��svE��<Q�w7q��zM쐗�q��N��/������˖'�.ڧ�M���s�=W������.(�¹���z���#J�E�ח=A��g��3��Ｃ,=��r���'�<Uf�N��Dψ(��1>L�Z�����W�7<�4�8�3o~-VD�JG{�����	�z�aϱ��c�i~��_�B9锥���#���P]=��%�^�:�`(�rR�s9��;ж��p��:6;�f�~��:TXR��$�^W]a�ёf�e��)���ꪲa�Eu�y��G��r�}������!c���v�"�����G�)�!�0f�Bo:�M=�Y*���~�op���~������.,�7W�,�ա*�%�ӡ�B�Ƒ�À�0�޶��z��r^����z��f��S�}���])/ ,XpB}v�=�Qx��9���J	�v�7A�!��e>�%󱆺$��k�U,�>� "d*|s��`�Ү�Y��P,M���׷�~��]�.����������VC}s�":FD�������%՘［�lyzk�������ʼ���������V����?P.�bc8���q������g�}�����X�����r��Ee�[o��1/�����xb��W^z�;���W�I�ߒ������7�t��c����Sጮج�N�ǉ8N���pĒӎ[d
�ᎇJz�5?�S:����.}����`��?�߲��/�#�C��������=�q���6�ʀ��Gy�y� ��͛7�Ҷ9�ҹ�����8����q #(Sg\g\�h�6��a&cm�P�.���Vg�p����	�N�F�=^���挌4�eD2�]s�r�c،R�ٖ3�s <�R���QFK�4.<mx���+Kg�#�t���逶9�R"R����D��a�!-�#@F*<I�]4?�9@\�L=�:��G;k:�:#n�r
������/b3�u9�0��ك�����Xz'���(y�O'�Q�V.]��~:R�逶��t@Fd���A�q�2�b(�Yʵ��k�F�@��L�΂k��gīKC��!���a��s�t@�>���P`,Jp�0�X'�^R˞ ���u�I�s�����}�K�[ �qO���>�M�J���c��m=�L'P�S�O~~��0�y0 �^�Fd��p���������ڢ�Ü{4�k��.�C�ĝ����W_�C�#��B���怰���ަl���ګ5��_�`aÝ9a}�-1\���se/�f����۞��j�)��F��<��ob׽-6q�UZ�fw֓�;v��[�^Cu����a��z��i�5U:ND@�M���	|bw4E�ВnOy�x}�\���l۶�֛�Y~}Ə�<��C�����N�[����K�7z��s���^�#�#^V�2�=�\����h˜!�sx1\0�{�G�iӦ:d�z������9AD3$c;0��	V�U��@��у)���b��Yä����ǵ3"j���<��@n��1�������%Ff�뮻�:A�\K��ı��7��9l�S��ɝ3r��Ж��|,����cN����#s�	^�d\�)z��`�T�e`��g� ���ҹʓ.Nl�T��(�0�+�� '�"�.��	�����Ç�A��^J`,��y t�Y���<_�u��7�W,V=����h�p�wXvڊ�h�1�m:/��kΫ��O諎�W���J3WZNa�2=���^�t�M7�c���YW�S���ٳ'~j�2�N��|߾�-8͜м�W1��`����m^l��]^4;;�Q4�s��=B��y�āG�y��B�=�7o^Ҷ�T����C2��m���9�P�Q��I��f@���+"G��]�uS��5u޽��{������	@�P<9��3�mp��P�{{��0ጀgL/L8#���9����#���y�8�31L5'y30-���L�3���LL8#6X� )�R���h?��؆��L��)���ˆ�#r�6�[;�ϱ�8���:��3�|������s�y>�z�����θ���	G��[1����7#Q��^���ʪ3��u��~���1b5oJ�@{��S}}}���k�}��՚���Z��;�׃���"=~�7����	g�s�9gsoo���g����?._��?8?�:��6mڰa�7�,Y�b��9"iܿbŊ�o}둱��R��Cq.�`    IEND�B`�PK   ���X���8  8  /   images/c52c1984-b936-4e70-81fd-2ef40f9d3319.png8�ǉPNG

   IHDR   d   ]   S��1   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  7�IDATx��}|յ�f��z���^dw�1�tB%�����	�� �A���H-���nl�ޛ$�Ye�U_m/�sgf�ve˅������7���[�9��{ǈE���K��ߚJח�:��it��e��/c)!����K�*�^�k����K`VV\��@!҅o"��:]��u�Q2���eI��Ŀ%H��������UTzV�a�����y�d��L�{���� B�%�����7���O躓acD��8��B�85�v��2���ۇ���^|��^w0ˇD����.Ѡ�(�o@�@D0
{�����3�1�<�V��(�z�X���ms���� �\M�������V��/z��K�"Őa��I��U�Tf⎫��������ƺ>��͉`(�L��+s��*`1*��;Mxty��0$��<h�GBm��ك8���vW��j��%��f��NĿ�WC���������l2��(�<w�f��w>�M�6�b������tE����X2��!���=�\W�w�����އ<\��������
|!�����_.E�Z���zI%�~p��d6�[��q��\6��8�"����R7Y]-���`��l<�����n��vt���8[J�"G%�i�❕�8&��N���N�O��y������\�FH�F�
�)]?�z*n�d���v��Umȯ
��TƦ��P0Kr#u�@�~��}�p��g�_�����뉍1R��l�K�Z��Jb���3*⣃����D[��D���RO�!�*:���FƢ�|,�ŉxbU^�}�U��N�B�!�h�Y��J�����_މ7ל��߰ eyV���w��j����W��^:w2��:�F���3M`��A�`����K�Pg^buI$�<jr����;t^�mN���tz�	`$ya��$�����b^�K|8BH�ф#�a�ѽ~OQb1�3�Xɠ��L ���Ѹ�AmH�d�yܐA�T���9����޴��l!�@2=J0���)�F=#;}�@��϶Eq��flh���w�_���>?��v3�}�I��"�ֵ��� �֌���ߨŷݨ"�|����Q���M���^k5v��m�II����J����6�W���'��[�
��*��]�%m���u�E����,�4��/�����N\��TP��A���P�m���h�����598����S�����D	���@�Bv���=��P]���ۛ\ض�m|����n dpw��E���g����	�W݌�v�(&��=z[4b(g���|����������N���ϩ��!l[|�)�?����7��׹Z��E���_2"��j���V 5��'����h��4��"�_�҄'^[�y.<�+�t�4��=��MOB�e(�6W�e��YUa��vr&��Z2V#&��q��<��PJ˼{ �Ӊ]�f��"�uʴ<T�"��"
Z����8t�Y��O)��l���Wp�5��
�'��$-'�l|b�O�eN�E���9��_�Hya�j���Z(M_�s6H�1B.���(/um��,3��j�Rj��V�j�M?~X��_܊��3�l��4��Hr��9���{���y���5X��S �6�M]�3e�W_�Sg䣳��
�P��x��4�����L��?�b����MH�i��8?���� 2I��tw�j�3F�9��S+����`�<w"��Lp�����]w�G~����m	��$�"�cd=���,����l�_v�0+�]>���!g1�-�]�&RmY�b�E��=C����������~%�?����	�P��~��]K�-�Y4�7���7�>%�>�<�`���(� ɛ7?s���"��Ѫ��b6�"`;�Xw�ᄚl��!@Tk%5��X�����@��^�<�i��x�����d@-�����g[�a5�q�ͿMz��<����:�4M��aJ��X������`~� ����̫�,F�T^
l�m��CUF�`%tk�Xի2�{7����H,?���C7����{VV������Z=A�N� �Z�R��:�lw��M�	��Ğiwz��T����e���+Z�<��Bs˰D��9?㢕A�
�q�#i����7�JuHƼj��w�s�s��Ӭ.!y<��|>����GhA�@��:o��	?��C�k7!��(��������0��,�Łu�"%�]C��į)��u_�υ��s��y����<�.����3"n��ֹΟ-��D��aX���X2�H'�<F���b" �doWT�ѷ��W�U-U��]��+V	���/�F���u`a�]�ɪ���!(O��#D�S����
RT*Q?G����3BM�R�+jۆ��g��x.<'cܳ�9�4~y����������bØU�a���=U��?�!�a%�d~/|�q�%�������;9jG�3�-��3ny���Y$`Yk��Вg��%^?�́>�mr��&j�>ReYc�	�F����)�p��A���t�
��e��*�%k9@��&5���YFg�Y���VebO�0<�cG
=�s�9�ܠڰ&�E���'?�ͨ�����[sceK����/d{	��V{��h�ۆ1u\�ܒ�9�kCr,�ZRu7����e����~Rd�g�=���Gq���� �n:�Xي�������o�L����q�Ǔ�P}A��ϟ��)8w���h��/����U�x�;����8��/ª�$s�ҮZR��%v����bq��Kf���q̅��@���K\>�o+KI����Ų�oŽ��*���C�T�́Z�-���,��!�Ÿ�Q���=���q�}���Uc_�%u�����o�#��!n�A�B�p�14�Ƒo7���N;��T�Sg����>,�9������j+/Y�xE�5F	����������_��S�Bf����+8VA�YhYS	q;��Ȇ1�6��	9�oB���LL��x\�+�A�s*(��sx+�2C��H�|$(˽��[�����I�>J�E%Rl��Ȱen�N��?)O����*B <�h$�	gb�k/fy�_��g��O�I��o w�,�\����,�W��vW�c�d��5�e���dd�J��2�,�^wH����aG�`Ua��}� �{�_9�m5���il�0mtz
�c�d��a,_߅^<^�v�y��~��֗N*ţ�q<
�<���/L�Sϕ���dF6c�����$ـ�~���A�_d�
�$D��$��`x-���S��;C��a�fO_L�Q�!��'�G�<��^>��5�6�hP@�'Ê�����E��(�8�^rl�*!d<J�/����!�-��3r���q�IQ-�.�P[�?���ͻz����@���V�委�����ϫ
&�XQ��yP�\�I%�_��}���.����G�(B,�/���x�#x�CK�g����.L��1�^����@�o��#�E1�XVlw��n d<��d&}�9O_?�`^��W%�BD1���h�WϨķ.;Ͽڏkf��J�Y�y��q5iϓ��� 顫���biW���&C]n��X��ݱ�R�f�KzG� ��q;c��jLd!�M�[��j�K�^?����,�Y[�o��(�U���e��
�B���B�}��f����v�b�䚩�in���"\qg�,kQB��d��d�,&�<OS}��n���J�W����3��{&��}�HU�C���f^��f���T��/o{�O&��f*�Glo�>"BP�t཮�x��s��@/�!�#��Q $V�&-Y���QqOאt���)⁝���HH9TwGWhN����������$,-�H,~�d�\L��#��#CB���ܣ�k��uSq�9���8�'��=�II��AҊκ}��b�U^�����;1�����t����%�b]g9���H�p�C[� 7�;'���?��Eߕ���{l�j����FT?^E�\�����94�/��?�bˮ�8��Y~A�a�»�k�gZ#���o���6�u�Z��%sr� 5�*�'�e�͟����W� ����w��c���yc!�lc>*+���'aNM������*U��*ad;<���QuE!���З���0��n_��[l�Ĝ�ōju�)�n���l����2��I3hQ�Z��AS�c+�RS�`H��EhLW߷�A
���ۚ����is�^uAb��,d�㜥�p�)�xk�v#�I������O��k�n��y�� ����4���Д�$��yx��N|��p���%}H��7-����)V�=#Sk�@CC^~�D�sP�Q��@E` _��+�8q�����~A��9]C4Y�d�m�~��"�&�� f��=��!>�B�����0Ϋn��f��� ����fB.���)��ǈ}��i��\"�K��q}��wy���I}�&eD"X���ܵ���S� ZZ��Y ҵ�T��9�:�P�@y���֚���#B�����ʛe�Ea�,4�E����T�~���3~gg_6�P��h�߆�`�X)Q-)��z�`5����y'�(;n������4X�z7��v�.=߹�J4�]��}��;���#-��h�N���zz/�&-���.�,BD�d`{�_x�=d�
{�|�H��):&�H��0��OI���Nƈ�4�sFQ*X
GeA݉�h�ߘ�=ΞX4�H��#ds=o&���I��}!U1�GDr�d̠�3D����[�W%^W �$I�����k;��"DO�ѭ�$�����u�&��g�V��v&ɱqH�L���N$𒔍��3�IZZ�{K�fZ�����,K)�pH41�� ��pX3��$�Y����m�:���h�y��K�Za3�:$.��Y���5�FK�Z�c�<QO�g����Ae6��R^"i����:��Mu������N\5m�p����;4gs=6v��+X,�����؉��I�ge����� �N���iX�^N��E![�=�ٟe�F�iAD|�S������4��y�0����AH� ���}�t�!h�]��@E�U������.Bי[ԍ���EnBbQ���)vs�C!D�,� �`����/D������*L0�b�� 9�=��ӿ�I��೏�A��V�*lSٞZx0,H�(�v�;�J�@U�}��e�QJ���7���=��F�hxI	����J�DHU�D�+?�D"���h"
��K�Y��D���QZ5~��6�~Z]-�`��b�i(�����>y��.a���`���ob6z�)�~:�	���Xŧ��4�0���^ER��&��u������Mz
���}S�&䏼y�
�i���*D�7OT-�����O}�>]Gm�Q��uAc�O������k�aִB4`[O�ICr�qRI+��ؽ�tw��b�1u�J\r�K��DD6���qG�z���Oa����5��r
6?&�uEN��d�ie���oe�&=���y2Ti��ٕ�is	uD=�͸�X�jtM���j~!|���4�-���Y����~��C򮜮Jє_�Dv#{�Ep�l2�b�Ъ2�U2�0�:9vIRW��~��j�p�L+O�23�p��J���\m*"�b0�ڰ���S`u|��(Z^�B�K#����g�LGC_^Lް��E%�ϫ����MO�B����mCY�;xP ���ԛ1j=��x膹�[׀u�G�+����� :�����U����akbeo'6n�GoO�����޴d3=~חq��k������C0j�!�J/!�0e(c@���?�H��DQS�͇��!X�������^�cf<y�	BM]4%-./�xrݨJ�(�E��HR��ҡ�(�
�ُ7v6�n_S,`���In�k����5o�h'��kgS��(� ��0�6��~��x�/�k ��}�"�t��2�2��2�������"Y8D@���sYꍳI�Uo/ס!� ���W�$��N*�R��r���&�E�ɠ��GQ@ ��H�cw�Cp|}�$��XI��#Ac��lq��[\���j��-�8W���<��E����3���b�d�d��"�*���Dl Djo�ϋ�7_G��}�t�;��KD�r�'+Z�g/676�=�%�&�6T��"c�̥0Z��L��s/����<L����n�WNy���T�;�:W,���n��v]�204�ܼ||�w��vgϨ���V8q�`Qe� H�I�	S�!��$����%j��U�m�E��!)��F�4�f�a���Ú��d{D�{r����x�]V9#(2��b*��$���H�C��#zxoS7��أj'��\N��h�&x��6l�؉�����ڣ9�ܯ�g'���h��)��pA��!�:��12��,Aq�0����Y4���P"k=�L���������������D݆�qH-�ءivr��̂,�~�Y���V�=v28��p�t,��r�
����F�/��vb:���Ѩ�:3뛞�	s�>E]�:�-.�;����R�?%c�����_��
V5�O�ϥz'��8���B���:��p@FK{��pR~��9e��}�R�<���v&�\����_�d��xv�f�}��8#�C|�x������O�5ԭ���U�H	�FI��EO�3��R�	�P�1#�j��ߏ����H��K���&׃~����Xꉓ�ڐ��|�Ϳ�y��K���$�fΠ�-�;c{o��X�MF�P���J�}Q�Q�j����-�}�x�T�x�o�[B�y��fL�Vc�+�@`�w�����%��P7EIk����M��;n4�p�-�k�L""&��z�{-���Qă���bdr�Q�e���@jaNA��d~&I��=�Ղ��� 2?���HBnb{N�]ݹE�Y��	�r���4��H���h�G��F,��|~)D�����P)ř�
q¬i�A2ex^u����2�jT4�kX	a���*`1UZZ�#dg[�,�h_�8��-�a"�^t��q�g(�t�
[̯����6M��9��PU��b.5J*�0�.%+G̾z��BO5+�T�=�\!�]=V�G[���������-.5�*BbP����+� `7����~������,X�yn��,;�!l^�"�#fNru��6�To/��31+�����Ӫp��U"5�O�7Zд�]�X�I���?���;��Y���y#B)���f�v����]�I�av��n~��H��TP��a����hv�4�I�����\��z�����)	�/�9�7��b��U�E�\��ښ,,��\��7�ioª������ ��چ�^In�T�����b�޶H���b���~�jF�5���*���df+07���H�{���#s6�0D!%���1���̦}�Ѹ�����'p�=J�6��ex��nKx2���gt�T7��ܿ]���	��b��\}�ۢR��VFE�)��7��&!wd]t���M�-��x]gR���:�4�%Na��*��%����(OY�$�]85{&���)�T^��$J�%8�}����}��B(�:̏���t� �.��Β�nvn�`��S� �6h�"!h�ͱ�����)f�ZTewA���>���0�����ErBr�*3���w虐��maj�����6c|Y|+IE�ҏ�л�sc�����J�5U�/�p��Q���ܽ��-�����.����A����6`E9*�c�1�n��^��O<>;��WC;���u 򸫲�b��|���L���n�q�e}N��16��sY5���.|���-2�/^X������������y����~k0L�������(r�&��(!�v�l%��-d1���!��Փ��o6��N����	��Qb�������O@�����qh��?�<`�������KW�}��aGAqdda���w�(i2?8�[3���ծ�/�]�\o���(,�J� v&�#�����Y��Y���I��!G>�ЄW4���M5�V�$��%�S�)��R�� %�1ruj]�-���T"(�����D��VOU���5���EL=un&�4��z�Ȣ�(KR̋�7���u"��#�XȢ�?�1E�i,=�"[��\ZeE���s�lBq�ԁ��D��r\�h4
�W!D�XH�SԐ����$�3e�n�
��QR1�)k��D���ml1u���q2"Y ��ȴ��}���2��(2����y}�YnCı8����oL˲8+���HJ�z_׊�&��N,�9��B�����]oo��~���Ɓs��h�'u�4�eWNEs�M-�ؑ���4?��M.�|�yn	Jr�ܳ�>q��Յ;��� p��](���~47�a���Ϝ{���}�V�[�Gte�aB˨�}�za�,g`����D�̭Oo��]y8F�v�������y�����v.F���[�D�c��}bnZ^��B�\6R��T�C6�F	�Ia�1G6�xV����)3
�l�_�ي5��Cw��$Ai^��j��J���x�(���٥���eكP(�7�xCݵ�8�k7Ҋ�2���!��u����ɠ��d7d ??_ �?C�"�. �q1X�{֠���$���YuEsL#I�����,���
ɱ�is(�/BzYu|��Ģ��	�ᄾ�vR�ƫ�>%2S��᫑�ă�¢��Z
�X^|�U���#��̛Ucf�\M1�Ė��G��݃.A!��4�)�C.���z��z"^ �)��x����aϩ��x_�!���#����^�8|BlB�Dq��`3�q�@EFGG���1�V��f�ɾ�4�������m=�h2�6��ͤ��u1ȪZ[͂�:�S�����W��p�b�A�}ؼ���k 0YP{0�Ŧ5���)�^ �{/���S��u���MAV�D�jq�~�t�#�]&�W���"�������~&�/]�˖-�)y��+�J�6�2`�dO���l��f�#�eĎ�Y�E����'��C��h�Ѥ{H����JP�T�R�%���~����٭��A�OF��Y�X#���mmm0�Lعs'�^/222RXk=��(���VF�!��HȔ���9���.}响��1��Շ��J��WM���ۄMћ��ߥ��g��!�"F�46c�Ǔ��9X�6�m������%N�.t	�=^'MnJ�s�c3g�Ē%K�w�^\z������x������.�܇�پ����G|��l�~"0���U�v��TUʱ��s���r+츌*2�����7��>����nx2�:`��N�6;K��5 �;}��,��#~�������4�
5V�`��������<�X4E��cm_�h;>b	r��,�$p'��e����m��&VFVVV
2t�x�Ød��Ԛ81��q����n?�>�����V#����v��ߍ�U5pd���֝�?P�����a���b�;o���ƶӄ�Ag�R���$Ss�p}hU�����B�Wȥ��1q6�Xf���h�¢�a،!��!5�+�{Y��3�Y��9�CJ�J`��!��%��V���"������@�H�E�},IHJ�b2�'O�Dy�F�I	� �S�MB8s��(���>z[>���m����R��"��>�g8�Վ���r�/7i��}��oޔ1�_!�+��,#�9Q�((������ ք�!��B�;�9ym� -�v�i�r��rv	=����֝$X\�(�3K�dk��f���@=��7�15��9sK���ԟ��=f^������{��P�w.�jm{u�`���B�aa���ֆ ] �+(TWNo�k�\`D��0���i�ɞ������?dL�A9*�',�hy�ULŤ����z�;1�Jj/Q{A1�T�,��)'� }pu�%U7߿A+iAy;ƅ{��K����"�'�u�S��kcV��U�]�EjEҲN>���}BNH�I��0u�L��3�ux��ӕֹ(i{&����&W�bC|���H$���^&"4ǀ�k�
�J6�Ny�Z�zԟ$�p8$�!Do���:���H$���r� �1���"e'�Q�pQdS���3���
	S�݊��"x�Am,c/�Jx�@iI٪n�x}�X��$��q����I��{�#�5L�C0H�mL1�ϫp��/]�̼	)v�g�o�i��%*|dE+V���i"Dٮ_fY�E�����Y1��G����4���5(���!��g��t��e��)�Q���S"b"�|��QX�za�x"��0+�?�F}�"\:����}p
d��r\���+9ksdIKI��C�I�K�bD�vB��Lm"\���+=�RnrZX�}ޤ��Ki�l�����v��1�D��OH�U���`���{��1�$z��e�@��*���yEa��n�H𓐲YL���2�a5�2�z��<�]H��$����<33I��q���Xؾʲ��i
�2����1�#tͤG�BE"�x[o+L\�H]w��nM�BX\ނ�,/���B>���j*>=+�����oiwP�~o����_�02N�h�e���!n�~j�L����ۿ�^��"���?b�R�]JZ�_"�ބ7�5v��O$wmc&�&m�UX�Eb��6Q��6�Õ�.�#��2�*tx�}��48��']A��4?i�Bґ������oE�
F�
ə��v^!/�� 0bO^����A��&��QI���|�gg_@��x��CQ��j����;����1���Jٽbe�O� ���1,�Ĩ)�8����#q3m&dٍ�� Y��e_Ԗn�1(12�Y��Y�!̙�#9��m<�TN�J𨒱�dv�8e�����`h%�Vq(�'46@�Rx>_:�T �OZ�މ���N�ZHs{{S�����E%���1L��uu`(hF�vz���]����2lFq�UY������1Hs�'q?������9�����(J�li����UY�T? ^	��eV�Dz)�Ԋ��q<���}�����$�4s���Q�)��0�ɕ-����_Y�MR,ަ�뇅���m8o��Ĝ)y�s�>�3kM$ğ�=C{�	,g_�75��y�X&&��� �
�x��,,ȘT�!~W�@k�7���!��q��q��|���$>�����	�XM@�q�,��;����y-?�&u��|4� ��3f��N��F�'���_>�L��+	�:߭�d!��T���B�pOo�`]�~�p��l�]{�M+���p!����Zh�[�T�Mѝ=��Ք�I:3���qYx��?K��.�@��@tA��qUxI��)*%�45��v� �h���ܸ�R1�n>o�,K�H#�W�cf�t�>�@�-��^U�R�|��wZb�H���Km�q��fq��
bœH\���N/\C���B���ŐM��Ғ�,b%|��g{]���X��U�a�1m������G�����#A�v\�_࢏�����A�$
U�b%t8i5<����T!��,D=)ڬ<��d�
��V(�����2^���"�r��;KH˃at#�h,��y%eĖ�
��>8�~�z;�iU�0��F�$���7t%�"B��'��������LD���_'XN��S���3=I]e ��8��i�<x>�|]G>�\1cѠ����Sk�pRY��y�H�Ml�3���t*1�51�O���3�pz�{-U�c:�V�x{�$�m|�~��U��D�a��b|��j~��$�؂�쐖G�Ľ͢?�|�4F��U7�يʬ!�,=�vL<yN:��ZD��j^��kw�]��)��w�x��O(tᑭsR�R�����s�鄣�5��aiNQ��k�*���_||�#D���I�d��7���$�[%9�]�{��������-4�e�l�Q�.�u�⊶̦�l|@T�2M@YB�ʓDnb�����*�|/�5�j2��27fx��J�|��Q�LO�"�c�3������U�L�@���ۖ�����E���4>C���)4��E6��N�AƟ�}�b���D�ك�F,���/�"�e�VG
����T�Q�~��L,���ɣ���QRꨍ:~Uƴ���qDq�S��;�ؗDuh|��;���>>��"���~�
����9<��1>���n�=u|cA�VVp2�.��3ߣ뢑9ϲ�&���@'B����w͆�7���U�Z�����=�B�ew�~9?���e�(���Y�v�|-�(nW=(MZA�e�g�G�E\'Q��������m>��q^���K�<����^�j�&��ep�vj$���Ue@j˶�O~Sz����~�{�Fn����ع��y�?�{Js�~J����g�o�W����ǯ��D��N��m����*��Q��  WKZL?�E~��3h�[vL��:>�Kn�w���E=�)����d}����DI�IQE�;�H��(4����W����g���5��R �#�ز���Af���U����74�/�}����>�7��Jld&��m'���S�3ǵ�L㛔�/�G�S=�I|�_z|���ٗ!P�)�X�	�V�w�|�K���,�C�U����[�%��`�%0�������[�!�୦��[�}gP;�H�����PI�̕5�3��H��n�A>��#��y�;h& -&Uֲ��X��G���ǗP�1BVѵ8�!a+ T,M��3��.h�v����)r<๼����4B=L��9�I��RX��3Pn$�0�e������͑z>��UT���X�i��g�o�V�����))6ſ������
]��/Ѩ�3���T'
S�kd�h¤��-~�=�{��X���.�4z7�c��Y��6���3�D�K|Fs_��&��Y�fx��ې���������W!|�қt]�7VGVh�abƢ�Q&�ۇy'�����C��7V-قm�=��0��_5t"�ꨞ����9�P�|�xhq����>��g�:lk85��0ϼ~ٳ�����Z�IIya$� ŃN�"gQ��ߨ5�����s��*����x��6��fۍ"%���Eea���p��#�u��[��	���^Wq8���Su��O�E���>aaT�:p���q~��l�����+�lf�x�6���]=��08*RF-����
�<������'�bS� ��B�x�ze��d������crۋyA���'��<�*�������7�m��9�i���Z���Cb�)�}�Ϯ��H[� ��W�=G̦�;pՒ
����{��t� �/��MG��\E�x�����Ɩ��F7��z��O�g ���h��f[D��M���4aqm	���]�4�Ms�ڿ�D`����B��(Fe�Ő.|C���ӹv��Ij��'N�o��N@����j>"��{f#PU�b� ��̱�*~��j<�z�@ /��iU�3��q8�x8J��[r�=��*3�[&��H`^�I����!��o?M�7�/�-� ��ر�u���N�l�m���ǖn|��qdHE���0�4@�as�c��z���❅�P$�dc*�p^Y�2Iv��
��<��.�0Q��!T�����1"��A�J~K'&p��u�׈w*2a̛�����ч�[#
�����qQ��*���DS�+�E�-t]B�(gt�B��B�B��3�e�z���������:��(�Up��|I�W��m�mq����(\��x�t��H����K~�h��eM�C���m���8ap�9E�P�)�{���D|�g�,Wo$�/~�ktM��R�Φk����K�`Y|�ST|�߮�H�&��z��-#���6�ǃO����q�V�@4}o����!&�n_��(3�4}vM�i���P=#������ ����NV    IEND�B`�PK   ���X$7h�!  �!  /   images/c6364832-c854-438f-b38b-75bf2a0cd33f.png�!މPNG

   IHDR   d   G   ����   	pHYs  �  ��+  !�IDATx��}	�g��UYwuuU�Q}��P��ò�[�c3> ��L�L0��%v �`� &�{�e�X�;,`X0�c{| �u_�:�Շ�w�}WV����է���f��������������T,��~*,���t�4]М�k}��%��n �-ȡ(�a 5n;*�t����I��p۬�4(�-\mPh �����	+�~'�oQPNľ�i�xcx���Ώo�ƽ]�hvP�i �BQ�vBI�M�O�os[��ǣG��Z��):���H�Wj1
�&�&y�G�P����
l�]�!��kjW�v�!⒥vVjg�/9j�c.;�S��8����������Z�!��Z�r�Cn���]�(�v)��dE�c$ wQ�e]C��p:�X&��ܟb���g�ѳg���ƪ=7�vp�"Yj�͛���4��2�ES��t���#�bzj�u�PU��F�q9�ZU�h8�d*���F
����6X�ǋɉq4��L&O��pX�V������ ��)d2��7 ��c��U���r	>&@e�譼�l��Oc��;����u���F���N��?3����&\nL��C�����!��#	����MG�[�J �ӓ�SZۺpr��H�?E]��e1�Jz��4�,X����n��>�~:��~�K�"���~�z��g�P��Fs��� �ɑ����,l���CMu���MN!�&�"��bdl���̂������ëZ1�A�u445#G�G�g(�NL"TgEU��D*���I�Q���(*�T���pvzfi:�]K�P�6��F��'\��kUĉ�����������D�����4�����>�������sb�b���ghc�&�2�[��_�gn_U�	�-����/�J`�e!s5�w/��6�MiW��������9��V�}E(Ni[o5�vˎ�R$���������Ϧˊ]{��,�S���'X�@M-��ד頾��m;wR3����]]�kE8HJw�|Xu��6L�2�����9��2.zf����ց���Ј&��I W^ú���zNim��Qơ��7�$��Q�Vw��K�x�+aH�/��D�ӊF�!��׃�-f�^�����6�0�
�Ȟ�T�i��b�#��]{����ؠ>�^ ��yltR:���������TN��Ͱ�%V�l������D}b�^ ��P�!E�?I��٭"<S9�G��4��Ժ�ই��E���*8cYN:_A�K8S���������	�T�@8����Z�FLq���fY������̣�e�,�8�����+e𙭝0�a�� Ǿ���*Ih��!b���΋VX�T-���܁�;3q�ܕȸ|�OC'�W�"@��\�7����8hGM����?u��c�L���at��X�ž�!��u蟎b8G[�_��|4��σ�j�ʹ�r׭n� ��DWc�^������Xa���&���i��n�h&b��������p��)2Y��n���(��0ZCU������R�St~(G�cS|t6V#20
�|-ɲ�&��޷wv��K'�\��-���/"569/Wu��yr��ܻ6`Cc-~�IK�tQ����a�������Q�`��8�?۹��n��p��ÉuV�omD�ߋ�Q���y1��� ��"i�A~�D��"���z�H��Ɉ氆��۸�p8���ؗ��@i!JRʖ A~������훘�1��EX&#H�r��
��9'�#�]K�3u��dV��M�B�U�d�tznT�gת:��;���_CX�;~����UȒ�fHz�^?Ԯ �������&���!	{�yZL��Ldɜ�p) K���5֒��[%3�����;G>�FDIҀM�SD��``��찘���!����vS������/s�� p�:Gj�'P�/�&�M��i7�nchb�f�@)G�Dc�Z$�ŋg����I�Tx�:X��3G��O���
4��&ȖO�T�J�w�ā�29�R�f!O���T��pD�3���H
llO��g���J����A�|��Y,��q�LG�$5AB½k	���e�>6!�E�p�(����Dd38�~�)������89|E>�%!a3�-1�+K2䏫S8�y`3����h0i�
=��*ND�񲽎.Ē%FL%��$�f0��y=�U:pa<%���'F��T����Q"3�0d`�/Αy1JQй���Re�G3��q��_��x#fHһPi��3׍��Hr/E��v��}�E�H_�}g�_��H4�
�7���^��&�7�/|�3�r:�����Q�mU�R���J7�F5|;��hO�8'.R�މ�t�U��6���cf�.�Fj=�'��
}�"CIg<���k��i��XZ8M��7�	|90_{�Y&�R��kT��X���cqS�8�`Ma���f��%F�)
�@b��͎��o&~���^��b}R)�~�����i3��[Ŗe�d�6{��2wŹ:?̜6aP�HD����Z����8�:�*�Đ� MQV�� =݃H�zd�������)�T��i���
���0m�n�m�ߪ�yE��ܰ��R��H����,6Al"��EÊ��!��33x���}g�Ŧ�}�!>����^��߿��`������f�q��9��@w���lz7]#g5s�����M&*�)�e13H*�>BG���)��ό\Y����m铲�L�M|�Z67L���c�3��i3���%0[��^[W����3����;���T����.m،qnB�1J݂����&Sf���.�A�b��� �HI��?,�q<�f�M��#�j���6F��$�	_�4�N���_&ЅXɳ%�d�&����KOh6�ia�3OJ>�$if|G<�t�%y�|�d��2��Y%fVy\r�	X�r�(0�����'�e�)K�+��Vg1��o��;RrZW��2ODy�3�¸!��
��Y��̌:��a
(�9�ϻף"�	��_<�,�;O�.�:,�;���={$�LPd��g��[��_O���ޛqφ�T����'��S�"���6Y�_�f�:��x�#V���9��
�6��O��i�_�TpqYy�J��gfwi)ib�T�n7��8�**)y�![�#����(��9�է��k����������ַ�k��6������|O~�����>�<N�Na1��o�h����I�vܷ�/�_ ).P�8�5uAѲ�(9�g�͉a���7v� �Ç����s��5A�����z{°��
�;N�G�+n��+2�W�,�y[�����6&��{_L�*k��g�p����?�߱A�;���Dߵ�_y�5��F�v9(b�r����V�{w�7�w<�OߺYL3�����%ʸ�.'��Ղ��g��˓��f(�v�QM�S�mg�r�;�S✍33Ù��y�1�Ḛ��������a>��w��|��Ib���~���q�??&����;�Dy�NSҹ}U�� 9?!�R����&�Vv�ϝ�~����!��5�)'%��p�n1W�f9�˄t���;���g��`&��.:XӾ�g�,��O`)e��&��9$-w�5b߹Q|���bj�8އJr�~:"�񼝋r	6�����lN��a|����>1�E�*���}��"�eq+O�q��eO�����T�t��4���@�L&�a''j��LL�w_;���s�H�ӽ�"�~/~��$0����>x�����ɡ�����o���i
8*ȇ���,��5�w��sz<�f�O�~6i��L~���)�oG�bKkz��1�|�Qr��n��l
�N;O_5��={:����	3"Q�kM67Ւs�P���ϒ�'v���i�E������I]f[9�������XC��~�%{��Ħ���������\�W�>�g��)\Of��������L���������DX�88`����Z��x��1ay"��hR��I��>�έ���-��()��ǑD@�ߤ)bc�V0�8�i:6ӱ���WOCs:��o��M�����H�9�KĲ���K�$>zC'�m�R�x� ��et�cPR�D؟���Na+K��<�~r��0�CZ��_�S=��]2M��C�(2�EI�����'�%�[]���5V��7J�������sp��Ϯ��m��ZC���FN�tƇ��G�Ã��g���׷��J������ꁫj����aUE[f�(7����Ȕ��(U��}�~�L�a���������x����)�1~��*]v�b6L�C��?8.����&�;ֵ���\6��'��j�y��(�0�Q���B�"_��,}���1�e��O�|����{���� �0-d�9�� �:�Y���DZ�ſ�;�H�\�����0�P���3�s��}�u;�r�whxS�Y�3s֞����	?�
�g1����3�f�,�2b3��9;�����\�(���KG9�\�)/�R�"�&���v�!��N&kϝ<�#S� x�-�cUx��,����|t��qe$͉K&
;y�����7��P�1TY����_��?�c'��O�V�U-�G�lUf�후1f��7�/;DժcY``���RT	c=�kJ77����?8���LV�M�Uʢ9lu�VL��U��*��('v���+��1c���1<�8@��a��t��m�5E��*j�+K3Ư/�����W�%��"�q��hּ^
{�뛜i_{��sU�R�S�g����ǥ�i�J(����� �,/e��V�S�����!�ݨ�o�
��Sc���4��{&�%�%�뫊�j�Y_�7`��0���~�"�.6X`
f�,�]�av���	��<��N�a)de��%�	]
l�U�N�4-U6Y�W�MNY(a{z�a4��OMƳM�e��_z@es��@!��@&P�8C���IWxkjq����_B�߉���D�u�^$�9�ۄp�*���s�h���ܗ�?0rA����ZWZ�H�"��3SQس)xm�+01�&�VDc�#�t��W)KGY�?Ȝ� ����(��0���ݕ�ȫ�u�|�~�"r��j6`K3Ģ(ט�� I�j�n����d��J>�`��n �B�������A��	ԫY���	/�>�E��7�`x`��Q�<U��VC��g��C�Hd4:~�\�Gjs�g^M�� ��5�����"'�[�y+G+�/P��J�!�xE�q�D���6 3%O�F�3�XW��32;���Sqb�&�W_c��<�hXuEJY,<����y�r�!o5pt��44��x�@�����]A���q�D<x�d�-`���ባg�/R�ѵʂ�>���C�ష��`������5��Mp�s�o�!�L'���(-��5X�)���~����S��*��?g��BqW �鋬����+b�;�w
�fL��czP��a�e(�p�4����h/Nf���K޲�w0���^��p��&��(��U�A�r�HF���D�S��	�v�9s��J3��wbP���cE�y�v��>�f��%*�	��"2bN��L�����hЋyٵ�!&8�S�nyg�$l�y�X�2s��_��*�*Ic�;��O5;PW�ď�
x9\���+�_^�E�3�ك�D߯|DKn��etD�:��j��~��3d�eAe���ɂT��J
�5�,��f�t^�7�sd9�ȥy���J٨��&;Bd�/`_�L�5�\6,�!���"��)��y�3)r\�A	(��ȼe9Hi���Ey�-�>D_��Wd�d�P�@�e╡�RIC��{.e�M֬�l�nW޲n�ˇ�����H(9����iooG?�<�_�#�5+%0ʢ�H��:��t�>��I(���//�'"&��TS����������*?.'�V-Hk���x}'5���y�T/k.]����֟;�h�.?R���^�9ӊ��ͱ�#��=pU+nڸN
�x���8���K���P)����E[[vw�¾�!�9݇�@��a�;�)���f�[,ڮw�z��
`U�Q��-�y��RE���̓�u����&pv?~����GQ][+�b��Ə~�#|㕽��l�06��g>�lٶ�͎O��G��K�����68�,���,ʐ�7"�H�)�סZ'��Hj^ۥ���V͙wfu��ަ
����B�q �PY]�O�٧����'�R��/��ؼ}�T��
1eˮ�x��
���p*PK���wf�)â9r�:::f�s8�L��D�Uu.*�#.2)���ҥ:�������e[��~���}����m؄M7�(eYg�#�͠���ݲ'��&C}���[,�� ��t%�K��`)��w�L;lW&_&��/$/�yn����aF3f3���5d��;;.Q+DGWW��=s��L+��1d����rŋ[0�0�b_	��)
-�z�p��5���bb��9߹�z���D
(3,�~������|��\�@�bL����R�*�%�xAx�	��}���r�̮�S���^8;,E�̂2����|ny�|(��]��(�Y�
����}��$:M������*:�8ݾ�-���a���Lb�G�Q9|���=s(���NI���G҈ݶ�c!Q3�4^�u./){x[3�Ul������q���9���2Q���Uu�g�9��p�����0���C��Ɍ�]���0Sjp,���r�j��H�pr�gNJ����]�]�MF�ۿ��fHYfCAY�u쟿�u|�k_C$���0JUB!��@���Y<���bt|�d��֥��v���B��ٚƛ;�LDG1���$t�E�/�]-XᔭmRN6�Ɛ�ʮ,���-.Zz�պx�i�D�P8.�)�����'�A��q�cޟ/����l���cH�"�C�_�iQ\s�vD�)�ȡONO#�����p��Ĥ�v5����O"�JK�v��6��Dcc#��uT�r~&6�&<K'K��|�Օr���XJɤ`��2�At���|�R�ᩞ��E X�yK�l�[��ZޟX,�JD.N0U� g�Lv򲉒efŽ��Ic����N��鸑��\1���7�����d\��l�_Y�x۶�KE�\Wᒍ@}���p���ۏ��fX[6H�SA���և�SIL��M� �]qU:~v�t+K��$Ō�ON�Z����i:j��睷�q;� :#'Vs��c�Ke���#�d.��ppi?.��1���
`�|L�4��?0S��vz�v�7�R���.r����?C3��&�sr�!��^u�L?.E�C���y"�b1OYj� M�ʾev$�5�%?1��q8���&�����3s��'F�?Ra��:�/�I5_)��G䊆<�,ȩ�OFxH�:k���YE�a$T�X��&d+?�`�Of1_�a���ʏW�$�� |\7���|H������h
Vs�o��B� ���H�^�ұ����z̳�2���j�*�l��A��O��X\�X��YԸR#�Ҙ���S)�x(fy�ym8
)8su���I��Ǣ\N#�b�p�5�>r~H�tr(��8~�"�t�s���#�%A�0�	25�|��'Ϝ�����Y�d�5$���z���35��p�!6̈́#L��S�BOdq�d�
u���ӲAǫ���IL�I}����ǩ˿�t!�T��l*�*��v؛:68[��31���	?A�}�D��s�B��B�{�i�m'�������B:����)\�!�N���#)U��G�@s}O��|.�Օ~1s�x�n��Nj���e�,2��}>��}7R��<�f�U�^����H}I%��x�bw ��I?��*%$ϤS訬㯠h����J&Q$f��6��u���?#�|��[�!�<dl}/�w���b!�a���zq���dR�kJYp���YImy(g!�ǎ�su%�NP8/���-[��_�9��[���If��`�#���Ν;)�Ȣ�p\w�u� SvapP"�M�6!FAƉǱm��9&�5}z|#��c���8z�� �i��_L$O;MG#��b玝b�O�<���fT�z00:�����m�d-_":ݯ�uw�!�������t��:� Y���w/�4����]	"�ljS�}�fю"����mb�y������ۥ�-�=ߴa���		�Ch�J��;�m�v����5�;I�,bf�>�ھMp�RKc��ċ�I�wn�j��֮�܅���ڶM�E��o�qԞ�����͍(^���23$)�?h~X�s�bb�?����#F�,��_.�ʸ��P�V�-E��U�|����/N��Q�C\�����W��)yk�����[�߽�9��h�@4����fJE��YDp�g�]��Sw���n�m�F����a��7!�3d�_揂q���޸~���M�I��)�G�2�_n���"S����,1��d%�³�����1� S���    IEND�B`�PK   ���XGJ���0  �0  /   images/cfd0a77b-9a45-4601-b836-f8aa27cd4ccb.png�0DωPNG

   IHDR   d   @   ���t   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  0HIDATx��}wxT����LI�7:BB��Q� H� �R��EE/"*�UAA�"(�{G\z/!����{/�:����) �w����<�����k���������������?��˟/kܦ��ׁ���
�k�T*=Q��^J�Dҟ����������?9;;��RSS(88�RRR������<99:Q��V������������L�ی��*�*����%��w~qB�ъ���ޞ��� ?�۫M��� �?|OiiiM�`� ###277���l�����-}}}��d��h����k<����rrrb�H%]�fiiI�������*qi��Ԕ���)//�)11��r9988PLL�|����%��<0F|�9����?ZA66֔�K��b̭�h挙���@���/��ߟ��:��������ׯ�Z��.��'���ɒl��
)�O��a�����c}��t����XXXP@@ �����ݸqC�dz��Mnnnt��uz��7iϞ=T^^ޠ�O�4����Gݻw�k�H[�`�ڵ�Dw�ܡ��x��
��������j� vvvt��mm[�70��]�
9s��50d����x�(���
<�2�@��T�r��mZ��]�iէ+?~��q��ϯ�� �Жnn߾=}��jڻ����і�۵�������>#	I����8;�yeg���=�i͚�iɒE��4��G\����l�� ��m�Vp�����LLL�ğ� VD׮~���MEe�Ν�����u�F��aM�c�� �w���q��dA�m����J�7���yx�^} QA��;"���B��O!�@�܏����Gff.��+}��:�?�,))i+��������՟��#;�[ HY^^�An^�n��J	7HI�5�07�omm��kG��ԉ���3k�m_���3ruq%#C(�\Y��{ǎ\��ߗ�c(''�A,}���ǏӀ�$��Bj6��6�w�6�~a����ڴ�t�dܻ{�FF�6t�ڵm�Z���IY^�c���g5!Ƶr�*:z�����*e<�#3�`���C%������-������TO�יC���_�ܹs��Xfq7�^F9_��� �����K���H�#�I���ҳ�x��.�6�|��UŖ��ȓbH��ԣGz����˻0/��lMo�9� ��=���n�j�F�T2Vєw�SG�r'X��\���"�d�1�+���&���M:v�EF�X)@xg���Q=��ʌJ�*�?Wӵ[!�9s��lm̨K;7b�ǽ�HzX�PIَ�vU�_���ѱi�Cy��k�:�
��Ҵ��֘�R9S*�;fiaBO�őB.c}g]*��~`<���XmNH�&CCC���={6�U��5dmD�#�t��ʪ��6�f�yE�6��v��{�h��ih�\/��xg���Z�0��_0�<��˕U��$�#��_���~��3������ʊ�����~�+�M�<���(#L����D�&�ꪚ��55w����,�;���6���|ц�C�$}�����&&�CgN2����G�6���bL�.���h?�����#}}�ၣ/��tS������?��������������HR���L^n� �ySS�cY�̘�q�)���o�2��������%s�<��"�<1A:p6[Ik-4&�#_
G6�>'C7k�����_P�IҢ�6���������`9��fdhл8)�Z��mӾ�+�+��¢����K���EU���Z�9x�EA9Y[�R��� �<�� Ӌ�ˢx�_j��D�Qɢ���x%��ח/�(�����@{;����m�O�S}z�gѨ�1��΢���roAA�K@��C4�؎��dS]PT6].�>d�1Q�6��>��R%1�og/S�j�&�����x��ӑ���W�[�iIO7���% ^_!�%+�jq�|����/������x�7���Ӳ�ս����D��@$�`J	A�R¬҈���{� �,G[����0�:0��q��Q����xu�ɸ�\�nǄbŮ�wӘB���3�i�B!���#W� �2���9�}�7vT��l{��x,,ފ���\�4,�rY�1�f�+^LS�W�c����c� ]��ՍI΢���@1�ZU:�Sq_Z�'�S���DX!��S�UܧU���I�ƓD���"�� ��&BH�20&.��}9�>�r�h��fN&gk���򯬬"C���y\����}_R�\�cu034����6.�s
)95�ڶvY�\�X�R����/,ՋO�mj!�I��f?MYZ~���1��]ޡ�	��=M`1�����i'��!&�o��%j�DǤ�/�4277���L���(g5F�.*(,m vR�r؇p��ǔ�H/656X��_,�O���UTTȌb\G��@2$ǿVO�U_�m�5�u��,��|+*�dhdN9�����ÇЯ7e��#w7�1,N��y���-��_s�?�����#�+��I���=�������[D{^��`nf<�'�`qB{]Ӷ�:p�ޛ=�����.�]�_P"ߵ�2��Ӷ;u�>��X�w��<lh�϶@�D�F�����+���L��5����ˏ�m� {]��N�6�0�笰��4�@|�������V+3�l��+B�j��(���v�̬���d?��u���#.�"�'$MJ*�q/G&^Y �{X\By�{�=��9>�f̘A�.��K��B!;�V��?6��U�}}����+���55Պ��J��F�.]j��*�.6���g�m�&��o~8����.�KHo@ D�/���cs� M�S������Q̑Vl�S\BF�6�F����C���HN��תǤ'c�F�D�g����L�9p��A[S�\~��8iǦe��F�M��nЏ=�{��*�9*�akO����Ix�;w�ɞ�L
<�����Ў����3�����M$�۾�@'���ݸIc&,�m�~�a��� r6$<�m ���W,B�U�`<�O^1&f����a���ذo�G�%�l�����護�ӥsR���;1N�WUWf<�Ґ2�*��TWܼE�L^J�7o]�l,�ĉ���I#�̣s�w�igj�ho5�m��x����E	)e4z�Bv��R`�9�.s��/&�J��ݝ��� ļ0���'<i�=ڀ΃7'������]����q�W���>-_�6��v�$�y��Q<�^�;9�.��K�������*�ҹ<�'dRR���MZB�Ν�˗/7?���Ǎiܸwh欅E�aTU��*��)�^�ק���v�����b�,͍�5q�n8e�V3r�(33�Z~]�R���"�$O�>�v��!�=b��"0��<yB�z�N$���(
�p�u�Ё:D�'Ocw��]�M+g����~�2�o��w߱4�LӦ-����x�� !��U_���E[�ncy�2r��q�x�?<��"�fff.�^^^ݸr�V~N�եީ��!3r�l-VH�����RP��,K&K3:|��^�>	<v�:�С��gݖ����w�Ӂ�h���h��u!V� �����dV����.���={
"Ȉ�հa�Dp��O�>"H�R�Օ��-�ό�<�Ol�X��w�ȑ��ߍ��B��lu^�z���Q�W�N�`B�$l���G��o'^�����gO
�[0��Wʆ��V�&�$%_�����'�z�12dqQ%,����Y�X	��1��יN����ĺʇ����H7�A����� �U��i������ԩSE��M"1v�"�����Ī9{�,�i�F�����6��V�&&g	�1�;(��)���<up $�,ݡ�zQ��h��~J�J�Z�Z
�@�QUT^K]xDg���Qԣ���h�/�+2r������OɫMw�9`&�,��<�z���8N�N�/~|���P~���Ξ=[� �8���-Z��8�����)''��=J�G�mo޼ɂDU7W�pP��kAl�]�������E���'D�իWY̕
���	pL뫳�Qɩ0?�������	o��E���mm^5�T�ʲ���M�N+�����d�J���əZ�nG	����ٳ��C����2g�2�=�5k`�J�nݺOQQqB$޸y�Bã(4��o߱� �o�.��
@<���T��B���Ņ?~�2�E�'�E����_~����|,���8j���������J����l6?~N.K�c�Iߴ�P� ���R��կj�����s��\�ܲ�h�B��th�F3&��jIR��E�����:����}����#��K�����h{�o$U�n��a.�d�"�\<[	���}��|GpmȳgB�@��322�o������o$����8�/^��,DTXqPQt�5z��� 0���md� �jZ�����B�O�"e��u�;uh߁��ӖA�ڵc'7�R��]��du+���R��Z���3U:�Rx�N�+@jΗ��ɯ���<�AOOJ���T�[�0j���[7�JA��|��H���.���w$BQ�ړ-#N��W��ʚlT6b������8���Ѱ���{��� 9�����ݭk�X�������ś���E�P�Ϋ��ϿֶW�YXX�¥�� ;�ҒC���8nUK���V�FӘ�������y�܃�(-��ZwC�.QԷ����L&�QTx�z~����BI#�Ә���i���0���B�|���9��:-��u��5�;���ŚNbٳ�c������b�U0p� �D\()�1��JA
�����U(b(USS3^��xM�x�l!E3���%,#K�:�#���HL:!�)suQ]^]$D[u�r
y|���J���p+��={���k�	1%���K���0������J��h�b�����o��� �J-�;'�_���_kA�q��"փ�"��"��8��(��XW�IEy�f>�~�5�3���ϛ�2ޙf͞O�~]h��h�I4x`�y�Ш��ћo��oѦͿQU�����K_H���WBǎ>ԪU�܉t1ƾ��y�	���`9M����<^XX��KQa�vu6�����H���pR7MA�j�L�}�A`68i� �����'MZ7'j�Q͇a� S���m�r3��S2iV�!"5{���V"%�h�Gn��H���k�bSH�9��w�o�j�G�.�f��c�C ��i��!,.���uXB�W�=�=/�D+�A'`�a��7����0B �+V�UW�Kc4^�j�b�z3��A���V��r{�P,Ul)��<u�>��{,z�$';[�wrd�TQIi�'��D�[��Ɛ���x/��{�A��
JH����峍�Ow����֙�[H��tR���}��	�PT�XZZ�W_}%<cM5	ػw�ѣ'[t��2e*[{OD9ӄ	�����l����!C)==�=�
��?l�/�r#�?����|�%�h��#x}�4��`�TU;��R�:E'<<y�yyV�dˉ��'
D4�?D�RT��5����4��1�_� ���������r֧�����
;��t���+������z*�NWݺN����W��oܬN�"`�)ƛ6m�0qa�UTT�O�6�Vuu��`]�W�Pnn��mA�O�8�Aj���+M|g0mڒ�"��ƏD����gM?��"�P[�G����H�r=H�Q!���1��{����։WS��J�/(fB���E��"�*ٗ� Oϓ�D�e98d��5���h�F�
���X�-����5k�"gG+r�\UZ�C����y�殙�!}��"a��cB�j����>f� !�~9��J�Vi`�Ν�1
�Q�o e�ΝT]��7T���<���,��"Hp/�s��9�蘒3��
�|��=D9,6�o�ԤH


���PXd<����b�@Ew��)&� )�(|��OkR%�j��㱝�TW{M���4#�a&D�f�����k��]���R ��;w��m ����/o"�6��˔����.�OWF.,u��j� P��g+���`q߫��f�%���N�e,�i���"���^����E��x�����%�.6��ڰ@�����ǷfQ����2(��n�mm����>�+ &k߾�D��mk�g_R�%�O�vVp5ع�h���`��<���W܃2�{L]��#��3��?u~C��/a/��5�&�ܼ����֭��x1X{�B�lb���ҡ��@Q'`̢x�{o��kk26��<��w�L���]������/A@�i��le廹�� ��V}ʾ���D"���T]�����׷=��F2g�PaQ���]\\E¿�	!�qqq�p ���5W �)s3#���� 2�Z���:���P\'-З��ueO��������T�:1_�UZB��%T,���5�a���1��g�i���<�%2��'�-�POkmeƃ7�Zc����M��W0�V�_�U�WV���`n�s�jaA��t��˗/����o�\�r�k�Ҿ/k�b58�j����ݻפ�U(��ֳ$�~^I�4� ��,��T��P�jw��;���r�=L�M��yGh��5"�6zIU[?�TUC-LX^&%Sc9J���7� ^V��0�S�ͯ1��4����(n�>EX�G�a"q�T�*'CE%�F$KO�<y^��J���P�f�HI)�	o��1!2Q��z�-^:Nv�Dߑ�ė��3��׮]����Z�E#���
�w�������zzz/��񮁁�5E���&�m�������,i��_��!���:e<͚1�.z�L�(66FD����I��}قQ��;�]�ec�����+�ŋ+�udlUUI�d�eCʯ�vORhbY�b���),[�`�R���ɶ";[sa���&Rjz� �K,�ןs$�Q^W��Ϊq������_x�
�։g/\�J�nܢ�g���FK�.e�Ċ԰�ucJjI�a����p���%$fh��k	�ܯ~ӂ\��Q��b9���~��7:�!k��ԓ�ESG���.�\!�8{u��:�z@���	����Ӹ5�3�&wQ%ٵK24�����h��Fw7;j��C�$H#�� :仟t�R���e���P#�D� ;��Bs��8��ݛ�)��bpvv!�"��UQ]Y.Lܛ�c�������~B<ܿ����<ȻUz�(�����@�:2*F�c�&j�P)��A���ڌQC}Q��Q������P�����<�C��ά=��5�w �1��0�&��+�.�!��5�"1�� a�zfeE�l�,��F0tb~[�_򅂨�Df��3ސJG�� �[������,��
a�޽��>D|�!�
����b-�<L�Ǎ��V��&NMqq�iէ�Г�A4a���>n�Of͚%B���b5����8t�����]���t�%ss3�hXS��>`��_��dem�]���]�x�N�<ŢNm��r��хҦ^��P��o��w�� �0e�1��&_H ~�k��ʱD�o���%�,8؟��!{�a��{&�5���H3��I�Jm��qԳ��(���~�����9!��j�!�M(+=Vę �e���J�U�[zJ���t���ΆU��|x~���&f�(9F膲�R:v�X����#����7de�F+>Y-8[�ԫ��X��M�-����iӦM�X���������{x)�'-e�==~EA��P��E���e�!fǫAr�h�a��n0v�Ș�"�<t(�$t�Pz��m�ԃɛ�O�[��ʪ,:q�i1}S�c,��t
rF�za1W(#5����Z�4.Um ����܃?�T�_�����X��=D6�x� �UC�9���-��q�}��R�>}�$̭<���`��� �[?��s<𕒜�,*~Z���3�"���}}K��e�@����&���#�TH!��P~y�n�HC��J�v+L�}��t�N8��"-���Z�S]a�駟
����̝:�.ba(��ի���ͦ��"�z��C}�4���֊��;�|�n�\��R=M�!��7]]�V�dee*����i��R�3+����|Y�:Z���K��7`޼yb�0��RnݺE7n���t1lc��*��2jĬp_�i�ݯd���p��A�bZ=����ݤ�`ST�#�}�da���JkàsS3K���C�9 \��਌��U}Ç�S7_/�jן�+dtj��T������L�C
#��k,��E���	Dn�{K�YهSzf�����oC�,j�K�x�t�WVH�}"� ���\�e˖�{�-0q�x��bF��x!���ϟO3g��Z�=��DQ!އh��۬$Q��TVR�:����EE)*E���	�U �@T/��rݷ�t��Ɏ�v�4�AW���
H%1j��3�z"����1���T׈h�Tn̦0�l��]M��������d�K���ۢ`Ϳ�7��{�����K��WJ����L5�0�Y�I�Q�)+-\D]_E�G$Nʏ�X�+��`  ����
�G{��jয়~5����"��"��֘��֟��5͜2;��଎��E���P����g
b�`l��(3�h�Ug;���H����HA挠YSzS+:t\�Tiހ��RI�f���6-�B���՗:�M��u��A`��׉)�<y��z�-�"##Eu#*��E�9V�������D��u�~��(�~���z���&�XHV��L��-�&���t)[���t!�έ��ܿ3]��T����|lUI�3+�D�x���,�ʄ�D��F�E`5,Y��.ͬ^�"C@b+ �	�g��/����"�vO�>􀨨(Q��z�ja������߀��|"(Ѥ�T����.MI�����JJ�>6�l3!6�T5r�a16Y����Ŋ��#I�S+�(>!b��-X= $2�  �G�[Xt�[<��TKB���l�@�0��o ��
��	��ŋE�C(�1`�p�ݻw�g�q��� |�ȑԽ[wQ���ϣ�S``�6l���?o=M.N6b.g���uqX �	lC�j��!��?��+ac��I�,��'��J),=M(uX�=�����|�8��T�Z��_Cܠbό;VLhv3a`�=���E7l� j�,�E{PP���w�R���O�1��oG���V���v�� %6c�,������0��N�*�M)�_��3l�y/��Pʎ`)5X%��zT\^!�|�/ؾ���-!�����@܏��}�6���1P�[&��wC,i"��'�=$�}���aQ!�@M�p8��O�:Mwn_����l�a<ԟ�Y�����2x)A�)�����-m��ۊdru�4=�=
�L3f�߼y3� �y�B�L!�[����0�8��<8������a�yXY�� � �Jb	_ &L�������:;v������^�ԡ�If��Sj
ʡ.��0O0�9h� ��ֽ{��s@�Ll�^�G*�j���ӓH���9Npu�1:s�W��3���s��DL��� �j�|���B-���z��(����zB_�?���;�M�6��/���;e��X�u�ˁ;iP��,��O�+�jy	�d�� Ow��n��'o�>����g�� �ԬY����-�,�#+��Q�n�f������'}��H@�v�gN���ޣ+���;qq�Mi�-f',��w�1����~-u��C��'] �V�-�o�Ɗ(**Eu]:�!'������)�I+K��A�յ-��!Z��B׶h���it��/4�O{b*���b���~dU��\���������H@��n�����(iҵW'A�A�q���j�Ⲳ���)lل�Y�3m�f���nߋ��"�y"S7]����DQc�Bcnf\�M�ع�uG ef���%��Dn.��Z��zق�=��sT4`h��y3ޤ.>�ؕ%��B���>-".%%�Ə�CCt�����0.v�hp4H�nmpp ���1a� �T�8pu�����h]��'y�%��.7p@!ڢ�B���+����b�L���%�1��
݃�@������54п�`#�b�ĩ.F'Ap X|\8���BQ�i#C����ShݚY�����68ZG9;Z?`�tr�y;>6����%q��:&F�G�K�V� �=v�;y`kͩB��Κ6����B���*��4�0s�Qk�ۯ=@�푽@�����Ue5��	��3����	���}[���UT�.)U�T�eC���kfV�����lm�i��� �!�*���sko��4�?՝����D�}Z\R>GkXY��8s���k��Z�8O�":�x:�����g�@Ki��jGk ��hoy���򢳣��0���&LۤxlC�����g'kZ��6m�~��~^���LUQ0�o+�����G�����*�JV���Tæ�z�!2p�	�g�Q�5#�>,"��'���#��ޓ�8��.]�}r��hMu-^|���Q��w���!H�yҶ��ڧa	�Q�;ut��!H�VNl������1'�7c���<�@"�igk!L�re�W�<H�T����MO7{ɳ����۟����UA�8�
�h������?,%I���'�����y8z�B}���x��$m������jV��c��(���'���2
w�����fNբ�F�N]�/v>9��S�xȁ��iv���Ĺ��=��?�{���a�����=�3fWn<3���(�!f����TD=���$��3���d�1�~�o29aK$��R$��R�:I�bC*C�u�䡋D[���ʣ���J�����Tezz����Zl���7lia�9���' =�Ic�:	S3�����dJN���p�����00��2MͲ�y$���� �5Je�1��|3#�Q�S�iB���`�3�eD޵�1�[TTf?�E��E�����nw��־�����ߐ�w^���cJˑ�����f<&��ʍ�"q@�Nn���./�4e������"y��^������\.jl��!3��~d<-��0C��Vn�l�iI����N�d@Z����	�T��k׮u���gQ�ÓԹ�� �Tc������%��VgĝP��Ȝ��7��u�;P�=5 f��gJo��n�Q�+7b��^p[of����B~�� ���  "B2��w^�:m�,�̨gi���WV����Mk+�7!Q����0�-����&h��j�V��k�b�m}�{�*ı����7P�SS�]e7n\��'Pt�9���
�x:�c8��ǻ(�زa�B�~q�Y�g��n�w�a������8|���5-��
V������ü�����>�C0Y��g$���/��EHDs��2�
�qwle�ɠ(�1@��>x����#�]T���Ƚ΄1�	"ɥ+��3!�"aA�oUꨪ����J^6& G436Hml����ΝO���b;����.Ɠ%���\��i�yƌ�����rr�HO�He��'s�>u�+���k������k`mm��An�/aqL,+�.��1�!Q4m�RqLlsPXTJ���x�xʊ�{��I�:}�1&x��~�/�����uv0��4�Ζ�
Ɠ8&���ԗ�$���)����X�Ÿ��8,���ln�8""��ڵ_�R>�b�q@p+c�V�E��&�����N�F_|�Z{f/2q[t��IDGa �� w�@gM�0�Kp\�������ksG5cq�� �A��@!�|$�4$"��q#�/B3����XT5~������ �8��6��6� e�)5��m�Дwߥ�+?A�Ռ�����I 7<�/���n�7o�t�w"�z��5niiKC�x	�xΜٔ��^�}1aķ�W�d09��[J�Ż �j�#�~�@<G��u ��⊺�I�}ԨQ�h � rA� b���4!������?��ll�Qrbe��Q,��h���`N�i��)�����fcY��~1��aٲ��������gxr���n�<tD]�Er�a�- AG��HD���7�2 � �t@�b�?^0�� X�ȏ����Ds_�/Y�X}?�	�y���ӛ��E�-����as��4��/�`����
^����F������Ba�܁�&�R@ ��R��R5�� �ʕ+�X��qX��=�|1v��k��m�g�U-��U�?�.�̞�    IEND�B`�PK   ���X��k�  n /   images/e6413bd2-a01a-4823-b22b-7acb31e08f91.png�{S]�m����9xp�'�kpww���[�����www���~��v��TM��ڵ�w�Z==�
r���>}B��)}�����gw8��OD�������%5�>}B��w}N�C!����C
$��u��ol�|�Qkx���,*���1<1�E�w�����8�
H#%PH�-0���h����AO�E>���1feEW���B���O�A�����f;��,��=oz�?[�̓����P�����8=�E
����aQL|��,�qƔ����z*X���N����{�ξY�p�蒈B��o�U�ЄK��:�HϺA��ޣ��G�*��r'9l\z<��X�)]X�*F��N��ѡͧq��&���E���5�d7��ƥ]+�8�`u뮟�m��2�e����@��\�u5¾����o�W����Ť�s�������z���2�3;����[ ��.��C�S29�y��X��h"��)���D�_�	��'���s�X�3��s�Tp��������@�?�u����K���C�۬ ffN��T�(H���e���|�;*�W��_P$�9��z�^�>��3�ZYvZ��tuF�r&��x�y�|Ěd`�~�,
[��J�yb�YVI�[��B���c�f�g�f3ԟq�"���)�hY�L[��EV�?o��v���ĉX�}�Zi�gsݪ��Zzs������(�O]��uV����v�h�y����uE�I�F[�H��!$٩ſk���c�؎:�`�h~�&$
��_q6��R	'K�-b.A%}[BcF��т�m���*߀�a��`���'���|X$3�+.�4;�?Ag���<M�SO��X�6�Ҳ�y��X
�.��z�N����o��}ѳ�'u�]|A��Ɵ��g#��mv���i��Mxp�x�Ӫ�b�bs<g4����J��~�� )��&?�u�!7�"��7A�#�gtt�P4��!)E.������7�Rf��YHO�mId1zk ��%0W*5�s����z�Y�q�C�A�e����Q�$��A�lۄ�>��T1nͱ�l��M�du�ߵ�J�S����J�{�T�߸�{�_
J�9������,(1Ρ1��s�8뤖����?�	���=�2�ؙv�R��4�!�azfsGK- �Y�"�Sx���Lq<�
t�R@��ʃ	���	��+4n��-�%��C��8	f�l�(�D��@�I�w
��d���C�1��
��(6V�B�P��� F�p�*>�[ �e������_�(X�����>�^b 7��H��IXzj�G_fD��Q�㇡��Bb�v(��|�y]|�K� ���U�Ru`̩�,�mz����A�h3��zPQ��p�o�m�PrEli%_�Ē�&��nD��#��E�e'`��G���S�`< �93+ʪ�|�~�adW��@��͋�cy�]�eR�p����Ӑ��W��-�^��V.fTy�v�:j�����ߍ6P���h�
?��qv��`g�&�6����T)��6�WaF�d�&C@���daN��^�:�3����ǯU	��GY��[Тe6g�,HA8�{-TmI`6~�¦f ���������&��Y��V�C�����eF���#���a��K��	))�������V{���k�b��d��9]rvT���u��D�`e�!Z�[a����A��?��'�un�'��v�����TƼߒ��8����M�4�*�@7 u��6_���i����?G�B�+�����;F�pJ���l@\`�sm �kgLL�`���̓���O6�ꮧё�Qdg�,�,ͥ����`�ޭ���~�Յ�6��f��i�/������U,�7Xu���9"�z�ÉtiY���'q-a6�)	z��3�k�1���O�������:|^#g=ry�[�I# ��7b*A.�u�&�d���k���'����⨳����fqvq	�l�RM��У�mP�97�B����"���㼲���ڮ�_��<�Y��u�_f�F?�y�դ/x�@�cW;�M�zy�6����KJ��$H��O@J�li��	�\��҂� ���53y3@}Vڀe����T��Y4�o�8-_�!�%6��,:"&���D���S��0�7n�(��djU�!�:i\��99C��(ooQ�q����މ����AE����37�r�$��Od������+F�:�<�����t!7 � ��}}PH<jT�+1�ɛS>��P��O��E�zn6P��Ӎ��HO}��'��+���'G���O�c�?+�v��?������o?D����Y=۟���;��}=p}#E�.�!/�֨H�l�5�r����p$w�{)���.�I�f-t�2�.Z*�7B
:B��^�l��DU0ȺlζJ��Rk��a���"Ve���~�偶]!�������c��OB=#�A�(�'��]/������$^8��8��0y�����nfna�bE��O���(T�2�LՖ;�ATVG�۪P�*�H?.���W��f�ܷ�$I\�?~�h����\c|��4�J����n������R�O�����rZ���~B��2� �$]ʴ��w_I#��:�ڂ5
#j�l�~���8ܨ!BT�]]����J�D �8��7!Ѧ�֣Z�Y�h�2�3n
1��=�=5�^�I�'BN|�nu���0��M`�[}��<`0G�g�{��`nJ^s=x�껷u������,��j>CG:j�ᯆ e�l�M��kB���!��c'HVҬ�#
�^�K���r�O7����-(7���y9o&@'D|X��ѫC""�3j*	8:i�$\������Z���
�@��9��d��h�Z��=����Қ�]���`Z ������ێ6�17v��։|�k#���͊��߯�9ًs�/�]�8%!��
/�@�|j��%t�a0L���f_���V�3Q�S}f P*�HE�xI���ߗ���a����?��h:���1��~F�g�E✹���R4�>f�^/�F�X ��Wֈ����Ũ���=�?9>�RѹW2[�}��{��W���Wn>;N��^7k�b��'�����D� a�r���'x�4��o҄�D��i�{2�|ST��V��@�#����B���t�4����^^�F"�����/<q�V>l�j�"��l��}��ӄ��ꆧ��4����<ak�-~VڳƧ{B?>�}�	K}��݉��Cy9mĎ�=��>���発��rdT�t'�:m@�y��V$6�/^i! n�8m��O����~X���S4�~��e���~�_ϖ\�a���L-�T�q��*�9p��k��`"�#l��雕�h�c�� �ї0��N��)��		�I�9��&���f8�ܿ�T;�Ֆ���KGB'qi��ޙ��0��8���ȣ�m~J6���W���#B"G��-�����h�j8x��»���&y�ЇǙ�]\W��^"}��t��bZ��.�V;R4�֏}�`g/S�^�8�n��$�v�·Et&>��z��&���W4�NS�U�Q�43�eF�l��a�5��ٍ�VҜ�x�������@���g�Ӯ^�:�"�z�m��.D��B�X�J,V"��*CXO���KH�|5n�5~���#	<�x��`q������SM����l�uZPo!:�b���}hѹ���Ys߾�D<Uq$�+<��#����2�V����a��m%y�8&YY�h-Y!�W�F�8R��le�TD�J�������E"�����#׏�TD7��%����z���e�]ϵhu��N�fL����h��>b|އ�RXC����k���XX�D�< �j!Hz�e]5��~�a�u�r����p���������,�g��kW�6��u�W��X�Y�������,�N�K���^��\�I�d�++1@�I*�lU�V).�B���r+�̣&�PQ����	3��8���K�h�L�O�)A`#%c����c�(:��RVnў��4����n���B�|��k���{9%���2ٽɺ}���b�W!0y�-��ܻ���]c�Ac�O/1�0f��:\��OF,�E��;1�F��!�}/j��6��a��H9w ���)U��〼��mkF��<%m�D�^���y8{�a��C�t����+�?p�u��ZS?\{b�;����!��%�)P �}��n@���2|��r��xGa	cb���W�5o�B�5sB(��{���;$����K�ѡ��	�T�xb�q'�մ�{!��?���N�B�Yj��ņd����Ί�Ε/�G�$����1w�0,���u��P���T���uJ�� �24\�&t�㭽���zo'�]]ՍC�xM�h��jA���m-ڦI�c۱���SK�F��`(���C�6Y�z9������N�^����l�8t����?P����|���w�����A �l��b��[�f���|���C��z�ٍ�
�*�y@<�o���}\�):�ٞ���&,��K�!^Z�hH��v��]��d�FW������W!L|�h?��EF/S��������X:J�^'
U�;籒��|�c��
gB"����R�T�;do]=�/9�dV:�!�ɹt~�6i��W��tp���8
Ӡ�S/dM�9�qT#����oeL  ��{���.$��tX�@�|E߉�x����X���?T9�D��P��(U�D�‹�ۆ�ρ-^�Z�N�����7t ��Z���7΍)ZL������彏��v��;�Z�N�K��QzI��?3X۶�������^۰z�E��/��Bk�xwI�V4ʷ������h�.gu*��#��	oNql[���w�t�VCAo��p F9SߤDF=N�9lDq�%�젱N���4GL%`�`T#9Z�E�'�m%�&(I>���M�����%�����s����G��Cy�z�4�v{%z໿�	h�����m!/	��N1l��Bs�6����E��"�DT:�`��7V�a!Nb�U�VF����i����w�����˦R�y8�F~���<3f��zsm����ZW�����RѺs\��k�G�&�� 9�Ÿ.�Gf�j����	��+��s/�ׂ�� ��/+�EȂ�1�8����1�P��(���+	����hb�� �� ��k}��!zk8BQ'��l�G�ո�i;A�۰*�~$���4b%~��<,=z�xsV�Ӎ)f�%耕]������n_�;�+�[�m�nl8��LT�w����^�K8���}K$�R_:�)+`���������۩�t�7\
��)r������Fڸ>�v�~\_&v?�f=駊��
�^�_�X����[\h�#����|@�Cc��a5�h`v}I��:�
�K�9o7<�<�݁��d��c���8gly����>�~��G��:�׃<�A/�T�^���ǜ*���}��������l|;�z�HO�B���N�F��ō�u�����N����q�w}�o�^~5��iGv�]A�/:�:khVh�����;�Cp ���ow�&s���ZV	uc~�o8�Ň����J�)��wܰ�>�f+�~�g8�q���L�[Y񍝳R�Z���*�1⥀�8�;s��)�?ز�l���*�
�"��dawj!��	��W��|"�������d�R���(|`]w�{M�����}��2�i{fM��w���l-�j�BF��5:<O7�w>2�������s׫�W^tC�'/ �}j���=5)GHF`\�0MT��F�L]V{�=�;�������~��JK)��c�c1V3�\��n.�����I��Ũ {�mm�I�uJ&=0z�<.>��c��kEo�zP�5X��i�V{,���M>�_�#�o��2�q�CPt}_j���+<8I���������?u�@]_�؄���V��#�f��K��ڋe�ZZ~�H��v�� ���2ck�#A�sm�^��(X�{���,3���j��E����K�m$ymS��Bw3E�7�w��,w��L7Z�ː%�G�<bT�P��p��� _�St����}]����Tv��:q�x�:"�.�ɕ���L�9�$";'�n�d��e,�����'�l���.-�����2EI���+� e;`�)W�~�ߙX���*�ն4E��[!w�w�������ef��~:J�\-ᖃ|�4����^0DZg��غ�U8f"M�%�j�FP3L���ec�]a)݂���_.�p8�94����=W�XT�'fv�4IG���*4�~ey�>����I��`b�D9�p���00v"��B�&D��"]D�.�'���#U�y��ܝ��Eeh�)|Q��J�����L'�u\��k��~�B3$ޅ��4بf�6����I�/��e��m�!
��}���jg=r��P�9�lh3F5:5�3W�pd�e����-ok�!�1�S+�W��}��aJ<��1�e�Q����H��qWty\}�Ҳ����x ���d���)�y;��0I����D��x" H����̈.��Ϸ��uUkI��s>�MF��x߰l��=��LMM=���|�K�Ϫ;��3��4���$��=��"_��ċ��Y@6��[���x6�0!{l�R��ѳvD����Vuh��F�vW���g�� OS���s�A;��5��#��|�M���t�������A�xJ�8/Pv>�W%����^P�~����A� ��Dp�����pt��O�o��^��n1:l��x/"t�G��&�{W�W�A��<�Nx���o�=1��!#�f�O�ϼ�|d�Y��-�aD�8c9kՆg�U�Kȋ����@@bf7��B���l3i�a������j������@�Y`����ːO°�M�C���̠�ηnq�z�C5����|�e��y�#��k�7�T<��C��L��Ijx�Q=�O���w%K�]GD-_��͇���m�&��y#Kⱨ���<�=�O����g$:>dpI\�cs���*t��u_0wF�]�E ����KUBwLC�;�-f6-�rA�;�	8��_�zx�P::*K�"�W��c�v�u�gkBЮ��x���_aP��?� ���?C �:m-�qܾ/��P�3i1�M����?#�ZI�d���=U2&<-d.n�j����y����/���{�Y�wT����^��j��
�L�58]�x3�!ḩ�
��������jq
�"�Y�6͂����r�Umǜe=�aٽHnt8���C�#b�p�~�d4��{*��3�E���Z�r�)��4�ypV�M'�!q��kx���aO�'^�'߂'b{��p���ur�F�Y�#��!f��dXwb�lWy������U?n���k&��Ӊ�~�����W_��?�@��S@�zd�ډ?X���oMc �$_a�Q�/qn.2B�Z�}Jւ\�CK�j���	�&�,����by�2)l�����>�8d/�<1nLaD&�^A��F��Q��4���iQR���1�&�W�x�t�� o�T�K��B������B|=�1X��[���<Úm����Щ3�5��ԃ�*���c������5o�ǩ��0���0���ok��V��#�}��8���qY����uñ�Zʪ�gN$dտ��[�si�P�߲��c	�H7V�
|^��wu�j+<�9���W��������:�ǜz.je�3'����̰�����Oo6�N���%�A���-Wo~�i����������)Yn�Yx�TJ��F��=l�1Ԫ51��x�{��mi���@��)�����t�58�eX��ͫO�I~�~;�+��L}������>A�(g��QQ4]�P����� 3拉�k?k�,�3���&$��p�M(�Ba,���X���&.Ħ���u��C���ή'o��ȐR�*(�/��������V�a8�ɢGχA����������X5r"ш�h7�f��([�������7��q���w�蹻�$φ���]�!]�~���y�w�N���|���2D��Cj��7��A0� ����A�۱ޛ���=��T$��w�̡i�3|8����5��Z�ܠ�D<*�I@#�׻��2)%��oÉ�K���>UM�P8BLrrN�2��#��pqAЄv��e 4"���Aع�u�C���cu�?�C�?.-��"���Л����0$<��Jpy��(�R"�B�w�N�b�I���zJ��w�=q�md�}O�1���C�;3&��s�oN*�'�@�1fU�U|�H'��>�������蝪��\�(3ƩJ��V3N"N#�R�J�>����,��L|iV��j<M�̋P�X�q+�[�>7fP��6�*qj���໩"�I���UåB��r�!�>@����������͈�j.��`�Z2���ŭr����&�wa��
1)'<����-��T��5�_�	�8��rT���,]��1��)|���ݺ���!���"x�Sfm�Ծ��Z+h��V�6��l���p�<�V��=����� S$�?,�|�JB`d�#f�-�������u{�Q_��/�|(5��ל����EE�|�hE�A�J����ݍ!����J��˼"���yk�x~���~*���J3�ڥ�h�ѣ����U���uc���p.D�Oke�gB'�"�C��	�?
 �q�ΓҌ�ڳY�l�w�-Pa��*2�ǓO �!��M����ɦ1fK��N�4�9/��ɓT�)� ��@��[=�_�p���kX�7o�3�Z��d����!R\��ӂk�p��)�D��:c)g�n^y"����Q��4:�jx�����Fl/�n��۶o{�������G.p��۱���;:��ݼ3Cx�&VY�34v��U����t��-4ҶT����f��QGq��}~�exdQ��.�0K|)B�'�LS,�h�V'���p��D{��"ߨ	c�J���A���C�)mZ��ff(�=.9oZvS�4��8����Nj���^ƠI(�N�L�r����g%�feOr�(݁˫�5
����;a�p��m�����ANZ������f���W�@�Ri&!�u�k�xBf5H�W�JOe�ھ_�j;�h2>^��AO%[934!�[���!����n$rDú����;u�bu�ߨώ�/���z�����g3����/�;��ׄ5��	d�"'�I��ȂאO���J*�@���&���{xFa<N�N�(�����7�̭
��КG[@V�S7L'�H���s�u��/K5���d�j�t)6}?1&|���+��'R�����5�'��R����C�7V��,O4>�'�*h��l9�w�)�۔��
r�{ʙ��M�e�	�=�-;kv���Xbu�a��ȑ~&,�M!���k�5	':
���9ƑD�߮QS���8r~��H�GN%$d�SP%��EE8��l�|X"/�:i���G���9�F0uy�5t׹uY�y�Jp�Dl]�w�����;n�����f��̬ I/�T��X����(���
���úb�`6_8
M�/�XR8̉8i�-|�\�hb�0'R�rHÎhA`.1�{����/_��Y_�q(m߉ěF��a�5���v��♒B-"�&�"P�=*e{�}L�o�R�
ﰑ��&֗�.�D6 ���ca?L�%o%%��;kY�Qki�z���k?*[�4R��ӥV�u�նu�x�w��i��y<Iө�//�Ժ�	�����ƿ�b�{Ȧ1f�)^��VšQ��-���;0�i�[,Ƽ�C�l"�2������񧞽�����Q	�K��h���\�k>��_�2��w[;�P}�<@=��&�`_�x��Ɨ>�	�zTA{Xh�$��ǯ�"��,�&!mX�T;3�J��&�YZt�kf�(+�Ҷ�O��^(i6r4J��^�P_{�	���>v�H(i�<%:"<�1�KC��ءF��̜%�D���^�L�h����b}i��95%5��~|��6��T�6ZV��7Rm2�M��UtH<�ȢȂ�(Q
�E|�<ds��BT�0�W0�SXm��$+S�~j���c/S,}��2�5�Y�8�c;��*vy>��E� f���6�y�F����Y\�M�J�t�}<N@&� ��>\Gs��[䴢�*�xj�J�y^*���ݍ���#4j�>�z��8nr��L�r�Z�+Ϭ�$R�-��el�p$�%���΋��s��L��癵$؝K�YK�A��$���-�œ5ŤU�1��� 8��Uz;�H	�`����A}��P��L�b˘t��{	�?l �E88Z��>ו��惜�X�\G�T��?���X��Y�)  *K������� �����v�C�B�	Y���R0�Tlu2���t��bM��R�<,Ձ~��/�$��1�UO��L	g*��1����¦ʢI�i-���/��Ma����b��jjk�w�a�7Pw�����Yl���>�0�2���ߨ���Gc�n� �}N��p���wؿ�)
���/5o6��u�,������s:���5vVi<�n�'@�'�?�4Q�h[b8�q�s��Ȓ���؝�Aw�e��4�ߔ���A�/��2\��ņ����9�������D؅�Cx]����$�n!��O��K8�L{$C�X���i�����R�HΗ1XM��	i����������%�����XYO��[��*��唾�>��G�l]�%�d���ǐ����	���(�Pp�_C\�U��2�W_��	'�+�^]픒(����̋o�b���4j������ϙYf�r�0j�̈�A%��8�|�.�0)D.���5q��ӗ��zW�����r)ɉ��:���Y����{;fnj��r[X~�9�<����q~���V�{�;ߚ_��/P���x�
��0+�	Hx���qE�g�[�y�Y I^�

IO�)��D$�� ������������l��De���tFe��д�� �r)Ӻ�%�"]�DK����D�E�Hג��(!G(K*���od�@:�ؙ�!l
��An�����J@�%�Q���<|v�O�r�%��r:ߺ���<p��J8��r*�f��nPRF�,�����B���1�X��5Ul�>��t���u�����Dr�1c��+:I������N`��˄SQRs�_*��4�"�5�&�~M��%��o0L<�W�o'S��f��+/�$_�NR38��u|c�U�3w�;�G?p��4�u����z�����w�%hT����8T�R����w��uh���$D���4��Z3{CA[h��@��T��lT�TJ�53F��OH��Rh%��\hp��ɛ����\h�H�~E�]Ɏ��Q*!�ouNN	�" �W�HS%x��.ĐA��;x.��MH��{3hU3��e����~�F\�~q��&��s?b���'ۄE��2uŋ���z���!�-i.�:�7ζ��<��w�xm��C���O��yu?�1�_\������4��s��v��a�N�����f�(�͘]�x���Ŕ�N�Z���HMAӸN�?����*�M2��b���pH`P"fO�nA	O�V���R��}�n��\h$ՠ�b$vEAGax��lz0Hh� �������7)b������B�J%lKQ�,�K���56ms��&hn�f0	�ŗ"_�����a�X�2�Ϭ�sD���|��z��Bb��Z�]�ȫ�D�zg�e�Z��!��[����%�+���N�"7⇒
����j�-���>>d��|��x���c����)��o����-9g$9D|'^cg����]�I��Z���I�9��I?9[©�>1�Gh7`F�К' �g�l�*��|�<�򎩲�*��9"�L3��;%�
��j��ՠ�9>��-P@ڦ��n�G��3��W���&N�~RCmuL��"��R(�J�% ��|!�j�񷄔��5"���������ƤzQ�'�o�-��;��*E̶v�g�^�3��[�Ơ�b�Ţ�.�j�����[)��K���4d?( �/�d��7T��S����׌�w~K�Ė)1����V����
8̫zy��������K�wL"�}_W��:�#��֊�Fֺ�H��?���ATd!i"a�A&ը�r�~N(m�0UI�-?��m�"�IA��_))BwɲLm�����_��I96ɔ�nػd,��2�B��͠i�K�sаǚ��=7rI�4;vbȖ�j���(��Vt�vd�O�Ն{צ%�C�`�(ȉ�ã�:o�rA�$�N����QqK/9b��r&2w�q�w`#Ow?������z�;�5�_�������h��8q����<�&s�N[����c�, 
_����-)�a�d��l�u�Eܶ34�����}Tb�W-���0z�[\?�M���3�E���-��9^�Z�~|�s"BBP����Lx�t}Y��z���r�����{�e�Pr�Qǩ��\0�c�A�-.�ե:��i���Jx��	3��<{~�b	�f����&_��uǸ�_+��9|�bjן_5�����Ͱq|�Z�3�9*�'kܖ^��v�§�J��'+�k"q���u1�K��Ē�Q����qK��r`�2k���k"��|��VUV�|��������?��������WHbK�൐7��>�[�,����P�J���~�קd����,�#��G���,��
z����h���O�{��.tƵB�'DGB��B3Ǘ��&_N�O߸�
�$�4�'՛�m�si�����(�GJ"�a�Ǖ���]��ƹ+
�?j/C���ɜ4��&���#��ٜD&~�=�D���=��)9��϶e�U�w�.�8-}�����Y�U��`��rl��홷��7~�Tj�N��18��'<>��a���ǉ�X������<������Q�ԮV&Ʈ%�N@�P֛�L@����fL�edhhL��8�rY��x�x#���붹�m����/������Ըn���|�4�
N�ߗ�\������h
�g�
�C�R��.�)��4����4q���(�֨-���c��c���LX�A��[ �������f-��3c�K�N}���L���	���-�l����b�����@�4�� �|;��$�"L
�y���������o_�)5�1�?Ip��,ݥ���A�f.rQ���D��HY9S��7V�̾S=���)t�5�Lh�;X�f�K��N���D���Q;�Kn��:zHRZ���M)ڎ[�R�MD� �k�j�C�'���\�˸�'(����C��5�M�5o��Pc��9r���w���;����,�Lz�;&��P�\�	����p��� ��� e��o����i7VJ̉��lH8�Y:�}ٲ�`�0-�Rs�
%�>C��H�ĉy�?�wV����V��ʌ3�BW> ���@vB�5}8=�u\�d�te#-�G�ɒ��s�t0���s�ۯ2�}���p0�Qg���F9��i��a����+g�U�bL��ݹ�c��ǯ�B��Zq��q�kʷ{VƮ[��fLE�a��A&"��� kIV.�P�P��
s�4������ޱ�xC�8�t�5+{�@���d�W�^%&�U?�S��l9������Y���D�ʂ���HG�����s�O1��]��,�{��ս%��cAADo���5W+�%���>�����-+W��a}�d'�O�j!�-Z�@(\<�R�K�f��u+�'��#��;��ZX&K.��H�ڹ\�f1��ߨ=�d��yK����*�ˇ����^��/�+?��c�'�Ť�#h��f�H��4'��9�uU/���|{Yn�
�J�d����b�h��*J,�����[��ڇ,�w���J�\�+�~?�&�w�A���,���-���H��ݶ����V߼�%Jw�K�:Pf���V�[Y�E�V�OO|v��H�R�FDw"��lb�/ )�س��S�gV�7t9vX�x;�p~���JZZx��9�k�;�Әݽs[��i����u�3�8�miZ�E�cP��iY��h}'��su�Q����M%G�y����ZwF�R��d�
�������R\*RQ{x��Y(E��-�+��a$�06Dy]H�7�pZTfM������0��� �L��Wz��y����kH�C�%"I�_DD�C�?�L�}~c��g$�5'�����h��%��,c����`�'V̼�����������:�^�F�Q�#���yezO��Y
Lc
]n��C�;J��³EYq��ʊ�?)ŴDTv�c���3�)��.;}�`���tp�)Ze8��v���:�5�y��ě��t�4�~?�H��{��p�� P�12�өd[�gP*=��SX%5�~ɦ�6�;"��cP�)~W��J\������v�c8>�&ٸ�Ѭ�f�����OL�|�9<'��N�:��h�8��|ܬ�뽌���Ll��78�u�*к��y�,:ζ�@ ǟ�Z�y��&�Q����.S�+�
yt�BDՔ���k��vz��>ܨg���h�O���P �uJ�y�ȄA����rF%���
����J��ߋ�q~K��td��m�b�ƌ��;�^�-��NWi��r�3�=���KB�yU�$!C�5�u�ϩ��0�IaF��s�,h���D����A�~T���X�ѩ���P��z��iq��ȡ�&⩉lv\��))�I	�G�qv�U`�-�p4��Y�����Ў�u���=�%�˻b���%7��3���΋��j%�^����_��eJ\�nK���\���q&w �~�&���{�ZT1�;m,'$��6�h�a�{��Z�)�yl�E��>w�S�y��Ȗ�f��IV6�C�H�3)�2dY*�o�Z{4Ge����{�*���W�g?10��X�X�eq��FT�Y�ߋ[��{&���UO�;}T�3X�e�L����p�gh�$M3����E��T%T��{T8�c��<��܋����<�ǔ l��R0J�u�28��e[l�j9_��K�t���X���%�IƬ�+�^��c�l�R�<?���Q��S�At���z.si$�����p�T�������pGhvV�=8k|�b����6O5��.�T�}�����F�P�M���-�)�Bna�ȳ,�Co26Г+}j���>��t��`PZ�\���5=V�!K�o��Z�w��DGg�xFn%��+���-����V�����둁���4���s&�o�UUAC5I�T�G���%B-�3A	����8�������0�UnæS&?�qE���E��}2ǘ�]��).�P�Pq�ld�s�ϋ��؍TЦ'�{�:�!}���.P8���}�q7����[)A�sپ�}q�7�0��3�뼮���;�q^�f�I7�����ˑORcCQ�b�`F�����n�D�;~ϐ��m��-
�[�W�*>V*�,��l�*�ePk����Zϙn�č =/	A�����o�����y4���`�ؤ%���Y��׿
��q˅tIB�_R�q�(�.�y �*� 8I������P�-+�'�(8�b��pX��.R�[JY�"M�޹D��:+̙��Ϩ��x�0�$y��`���;�vF���}|Hyu'S�L�1s$&d�ݏ��y)8]��a��&��(���D��4G���(L;2�o#��=���_����RJ|i�q�� �){m5M� �}���:�1�jݛ�=��:m@��\)%�07�΃����~?]h��\��4�?h�e��+"���bؼQ��9;(��X��Dp(�r�^�]�0i����W��3�⚸T�HO"l�GL����Hi�O�{��Tٵ]�����y�P�A9�?�$`[�P:Eh�<��(����9����	F��Z�Q��{�B19AB!r,���9>��\�K�����lʒ������!-�YD�����q8�N�49��@�g�{"m^���.y���������`��]i����j��]-VUM������l��ol-FU1ec��'L��ʉLW��rϬPxN���?!G�Ұ�M/^]�3�K�<�}Txd[�Q����۬_�7dB��]#�����9k�<Ǖ�R�����%�ydp`��d�Zᥐ�e���"V�u�$3+��p.������$�K.�R�&�N����S�S���}c��]A��f� ��*�`�0b���JV�9{Ǘ���{Έ����>��!8C�0$�˴�XSw�z'��1��2�&]��8e�a����|TV:r漪oE8�� �<hw��$b�*G̚FYZP����k���X	Ӵ�$�ccbLlsb۶m�ضm۶m;�X�ə�}���p��Z�ݵ`T�+e��y\�6d� a$#��Y�F�������m07W��ӓ���}r6$dD
韽[7��Y`d}mM���O�Gr"';.'��V�
�LK�,�i��@ 腧�)�tԣ�Q�5���7=����ǥ��&��
7G��5kZ3 ���Ro���S*.�F��&�F����E�蠵�H�P��Lg<`�Pd=�oM2�`ȹϴ�hJŖ��.+�X�����!�S���qok��Ġ��^B_�`�q�l�[�H���d���r��Q0�����^�mkiWB�`A�:O��T�A#��y9��*�0B�����Og$����*4=��EJԁ��Zg�j	��1���w�R�������u��܅o]~�����$����Z�|Lv�����q@�e�J���z�2*{���Fǂ�)�D&F�H�
�C}�Ic�3�}$�p_�_	 �x\�=�H�s�ۑ����n4T����t��hkܥ��N�!��-�r��%�x�)�#�^��a���/Y7�])E?$%pf�1�OJ{x�i���2�ހ`���ɮ[�� E�Z�rL��I�,�I	���>�oO��K��pI�����}\a�D��K�$����$'����$ �!AO����o𹉞�׾3Q"P��c5B|�VPg�����0��XQ��~����X�l�^�F��C�z\�n����< ��O6�-�{��{�ί�>:\��*�N�x,����%K��sg��K>'��`��ʽCE���i�}�V]��$���}�BU9��(I�բ!���g���a�������k¦UER��?����Z���c-<�k�,�ꡫ^��-v#�_U��uG�IY.���M�t���,yRys��r��p�|=[�%�R�׳�bv�P��z8z6�yz��e!lK��Cߨ5H���Ȕ�q�V�t������p�%N&g��&	U���"��=����w��I�v/�ՙѺ�c�dߏ]y^k]6; ���܌���[��?;��r^�rǆ^����hR�I��RE�g���qH�%��$J����ؒ �t�pn>r$r��[a����9cE� �Y�9�Ἕ��T����f7$e�>X�!��QS������ZI�x>y�e��-���$��x�$��)紤���_�#{�C#k�l�6�����a]�L�h�F��Jc3K�\ͅ7O��/,c��	V�0�;Ѳ�؝Op�B�x9����xjt�g����2���P[Uv�bC޼�uq�ɈBQ(�ݤ<D���k}77���	��E���;
����p�n	D�]�˨��Y|-1�
u���-�\�a��@O��;#g>^0~��������<-"�M���=��?S��ؕ��휔��:��|x���"[��{y)$�w�q�}h�`DN���������r�c��/_�Q����;/8ۜQc�5NΘ�B���5Y�ɋ��̈́A����/���K(FT
� ��6<	H%
��
�5yP��_Y���(mI�9�1�6ֆOC�l���̏/����?7r37\x�{˝
�(*��&2�l�5-qh�*��/g>�`^b�;�ݬ���,��=H'9_ԥ5��͌*�4�De�MGJ�M_�ɒ Ҵ[�zr!��:?}{PƏ��*�y��D�YP�$���\B,�*7�_V�T~�֯c���_���z�لf��t_�����7�z�x����:���M�}<W�Li����z� dTe���C����ѫ��'Ǥ6�@�����f�B�z>"���+��`t|*t�u�I$�es��yyB�M��t��c�*��=S�U�B�g�oښhP�Ի�����꽽��FiY�ɀ*kR��>*ߓ��DzF��B};^�����%����Q���ʡK������J��F�3���S{_�Z#1L���a��{�!��N�b�Q8a��5�CVR֒�L����"ۛ���f��TNFB�a-��������m�O:$����?s|��f
n���Y��e�8��B�	!j�jyx$�yۯN'/e��;��D��"�go�d�̇?�]�;Z�_U��Zz�]�'���;���v��h�����񌥆{�-�s�hnn]�K�D#f?^��:�z�J
�W��0���#�;�̷�����;R�%�F1���d���?��8G��U�������υI'�;��֝2��5?FXf�"ܵ[�@��t'đ���q��;=�ٍ�`����5�@�u$�&��PB&�oT�7fR����
�H�~>��2At�&�E}D+��Z�#uߚ��L�PAɜ���p32���.���s^�XJ�!�I���w�� JF�#;�R���t�=i����1����!_�	&d��|�#���^�[pݣR���%%x�Wc��?g%�!�q��y�Z�:r�R$6�J$�h^z���LF<*��	���֙���2vn�&��If�Ӿ���5�a�6gd�S�Br���|߁ӾÅ����2��b]����h3���UX��kp9zB�L���h�ֳ��m�M�S�����$�<���v�>u"����� �/��U��=�.7�� *!AV��
��;q��j�)M����dIh��&�%�����d��$8D�E�{��$�q��ݑ?,I�?!����=vK5'���d����>Y�a�t�$4&XȒy1�$d�[}D���f��=�zW��<*�H����+&%Jc�z�O6�k��g�o߼��(�#���L%눝D���q�;�1��3�G�	�������#�����ET���%Q��Ol�����q�8ٷ�C$YR�
dzo�P�q�L�l�\g)�n6T�V�J��[:;;c����fyA"����G�N�/~|�W�7�G����,��[ħN F�]:�;�)����_���v���k��m��!���x`G�y-n��ͳ�K�T@t��2�A�.�Ւ���Olm\؟��܁UfG�9���b�޹��S\Ǔl�~Կ�p�����=j�10ē�⪧ጵ*`� �bP�?ͤ�|z��� �1X����Ƽȅ��*�Z�X� {�+23�3P�?Y>�hX.�S�V��d-�������=Y��|;��3�,�d� �D��<�Dw��Y��:���:�ܔ��&�i�����V/�WUPK�%.�$ƗG8�4�ݓ��2FEA��[�7����O�D�����[F�H;�Ŝ�y��Y����7/��3�5�sP4�N�n���a�JR�M�'����/R���?b���O��>���/�������y�/��0CR{���y�+��g�c��r�qW��Dw������vYP��xށ7�7�Q��ǂQ�!|M��z�N��[eC�;f����*��s�z�'��\����\B{T\�7x������J��_+&'�H�v��"�HF����c�"���2o^���M��@�� 1���x���p�����������Nw8� DD��US�x4��p-�0��!����z#�\[��`�$�'1^�2��!����馲���.��g����z<�-�7�	���ٸ���A�1�
7��Zc=B��L�XR�8p�|-�M'p��ZtB�Z@����:�xؐB��x����ۃ��Z���O&�hο������:z"vl�lF���Ԧ��}��`��R�\J2+L�J��%[r�?%۩e!<Z$��]*	���]8�7��9M=�7e�vR���a#B��|����j��wp1��/]��B	�\����l��O�^ȑ�P�|{���M3��]������s��1Kg٭B�>��FoO��b1�ݮ<6�R������~�c{]eQ#���ms�U��a���y1"f�GKN�'�P�a�zDh�Uk T��h��
WxK�zY�3$	���1S(�6��%E�5x�������+�'Yy䌉���\�0�*��2+����(��5�?����3�U�w��6�� ��ꡲ���VC��F�U������NA�a��e���!���(0���)l�J�a�foͪ�ۏ	6+�)��"����.��%�!��[�8f}�X~h�)p;�@|��wBI�Uq�A8�!Or�*����L4��Q�G�Z;𡃑�������E{�����SX2[8�2���|�_ܝ�R>�Cՙ�BpVb��i�6S���G$���=M��N2��8���p�{�p:Sn�c��2e��@7�y��$2~�m��w����[��y���:
�כ��}�=�^߉h
�b,�|`�&��{������������;���w>�+;χ���M��4 Z�$)��4fOl�s!&��?"��=�KS�&W	�.�I Q�]�؟)��ZN���@�S�zFј�{�/�l���)�G�Xg��@V�0��'�_�x�"�'�4p�*B#Vy�O���<<v��P�M5�����k���?������R%��L���S I��+2lj�ң��a>��R2oXx|���_]a�YKط�u��Wq�]EA�Q�I� 	-lu-��=s)qL.���zV�E���I��=몮����z<}a�TTe+b��^�g��i��yl�¸I��zJ��L�}a&l��Nl���'/��ICN�R�X�]�2���ڡk�s�(����S�fu��0u��F�Ŕ�|
~���WM� e.�OϋD�����1�;�C���N���=����lb҅�����D�Bؗ�iD�׻��������-T��A��.����^CY`+Q1���rv�������k�5���H� ��r��w:�y��P�������/"|~��|u���rI���n,�Kz,���.�+H,�+7r8+V��JĐ��(�=,�Ș>U�;�<%��s"��mV�3�m����Ry|�� ��-B��ڕ����<Hj���ߧ�2��2��9��ꞽ[���lL�4�Z��
²����Z�Uj���>��Bӯ�^@�z�"�Z�񉂴I�:�e0����ء��RjX���Ì�?�8�P�E�P~8ͱd(��#�1I�yR�a[�W�^���ֽ\�ihX��$��k1��������/�Y�Is��t�-9�a�7u���GS��==KXØ��G��I�&^ν[�ɧSD6�'��w��	
�2��=`�2i�<[��m�$��Pj��t���n���0��H\V�Z{��g8,1[�V��L3��q#��2.��M�ƕ�Ñ軬���ҋa�;���Щ�j��o���"ٻ�~�y��p����4��ǍM����F����@%��:�ḌZ��	���7�O������&���25�����rh6��0�t�s���K��n�o6m�U�{��B��/��l���@)>]Zᕋ���X/��LC_�Q�C���w�(�ոR���5$�\�2��?H� O_
E[F�uBeJDF��U�_�+��1�4���A����/ ��wfM�e5����E�k��3�������xc#N� F�d�
��(qo8nL�%�/�q�':�t�,3�< �-�I�ڢXG"��p���U�rw�����Cc����0�4��3�s�wܫ9|
��T�i�1�&ư�+(��Pl�Y����)���a�1P�bt4�,˽c#$ϕ�׍	kPǨ ;�	`��A�_���1@'w�Q�>D%�u��L��% vY�!���7����0(<3�����O�H�w4��R������ʃ8��cy��b���N ��>yq��Y*�C*�,tP!S�)Qu�4]��C��!L��P�����SZ�R��: ��x��*�&dQt���rd G�����uA"dҳt- b�zR��U>k��Yz�D!2���F�.�l,x�;�L%(���~iol���淈M*��� ]����F1�P��6c�:,)vm���fɛԀQ¬X���b��Ws�S�T�n�t�;����H͍�5v�V�h������囃X�H����k�uL�p3�A�������qt����N᦭A���iw�c�����)��<7]��f,��VG=Q��+w�K���fAkh�cc������xlϱ{��q��'܈�"�~f��E�k������!� (�&�.�H�<'�sž����{�]W�sM��;�=׎��Z�$����?��ͩ��agy��bO�|>�x?7/�<���7���K���D�M���e�*m+Yd�I�(R�����W����NQ$�1 =��C���)�����hP%_Di'�q�8���1�.Re�E�^)@;`�3�P���ubd
 8�L렫n_.PW�*�f5@H�G����b�t�A�[���Ʈ2�(��E>��ʋ�E��SP?1�p�\��l�!�w�`�/a6o�'tM�Ω7
-�#�[��K�%�G�g�y���	�I���c��[���J ��l��ĵh�̈U��M@�K�"!q�E��6Y Dic�U<L!�{�Q��~���m�=x����m����jb8Pi$U�&���`�N��z���El�3g�ϸ�)R��R�q*�n8�����&���ۗL�����s�R������۫�gsϿ`}?�>���S#���F����N�Bi<�����)�� ]s���n*k@hI�8��7���w�m������X���q�����H��P�<�!�2����
N\���|���߷<���p#�u� ,�+���_7�zb��Dq2y~ 2�\��}F�p8��(�n��8���ģ+u��ܟ������.�􄠄�=�+�y'��]�G���d{\Pu{��ճ�j������a�٢�`R���6$�/.gf������)���k�?$V�k 4n�\l�^�_�����N�s��?�E���13��YH�Yy�������}1��@����0�ܲ��3��,�
�׋M�Ɠb&&���b�~��=����seú�x~�K11}��$��}�B�ϧpw�̗Dx@����F'�8�l�W&�� �H��K����G�m�e�� h��*��kG�u���~�� ��>��4r��J��^#����C`e�BC͡E�V���q��u�G������h`x�|���L�+5�hG�`��J����0�Y��f�������Ak0����~����z����B�Aq�>ʯ����I��Wr���@���Dy�b��j�z*��,�����g�N?e^`Z+Iq�|M�jmA�Ji�c��6l��MP��a�T�B��"+&`om%�·):��ԃ%����G�[�N<4n�N����Νe�骾mK$��j�g�(�U�|�����	)z�a�m
��qdS�}���c���j��I��^�����H��x������o3�X|5w�X��r0{�ǩ�K��L�'��;U�R� B�Lzڄ��K[��d�մ����|��G�$%�L��:_�a��:��8���惁5�V��d�{<�ބ:O$�/~�S����CT�xκi�����ß>=�Ǔ=1d�X2ɯ M�ձ�*a��n�4��&Y��i�T���)���*g�2x��e�;A��i���eۉU��<V�<�W�{Һm�jAm[p�>���3���㪿ّ*�nj�p�}�΢�j�4��0�ſ?�
�g
��4�ƒz�NڤE��
�ߟH�K7l� ,�����p|�0 �TDbnN�#�T���|m��k�?P~��!��υ?R�͵W�5��������b�"��n-:z����Yb��#�܉�����!��ZDRc?<���n$-�9�#Je큐����A@������3A$��D��NF.*�Gg��=|�>f
,4����v���\�	^�ZP[NQ?�
�#�%�fTΟs[�2By_ت2Yn�k?�b�[�����V��S짙kpv����.f�Qت{պ�8�)�I<��f{���%����d^�T*����:,6��>��]��N���1t{1������h��~��}�������_���8�&!�ҴעE�aT/�J�\ƽm�&�@`���w�C~�R!?,�z�攠L�g[��B������Ƌ�Lt��w1*9]�_u-YS��X��Їۘ��7h�p��`��b���t�����|��D	��leR����3H���6W��t�dR7�h� ~�͜�;�K.�R�A�NW�y}�i *�=�SlBf�h��S�*)�;��X���A��ڏ�T���V�d�0[�Ե�[�oPHD��������.�o�E|��Y>���<�w|~����D���yY�	W^`��w�qi��3���|~��.}\s����C=�����1�����P����N�3���c���O���F@I	�l�:��܌M��7q$�B���������q���5��~��^�z7�vP�m����BeH�['�2����T����cGL/j���>�bm�O�q�1�01��5Et I?�m�+Nek���T����id�dQ�#��m]CV�J�
�_~�#bH�G��OM����j�F���գ>�gS��>]���k�}h�@�<�5��~H�N�ξ����/�v���4�3����~��^�!���֐zo��{��.{6�n�c0Ig�>�3�H�(8�%Jlpw�e����,��P4`���hw^oeb��:[�����>�k���������O��^#�w%y�]4�3�3wP|T�?O��af���=�~!.�'൒�lk��%|A~��g,ڎ}o+Ǐ��B��j6m�<�����G��-�Au8v8�7�tW-�z?�7�-%����n@�/J��uXX��&������7�g�ט,�0E�y��8t�U�=3�������N���0��{�8�=�=��Z��9>��7�L�5p�;u�Y]����#��dE.�蠄�O�lL�Z�9ӄ0�q�/�}��/��r򯺺��n�yn7h#,�蝈G
rV�Ĕ�pt�m���Sγ`�b�`;�C���(N8	h�DF�)�$�~Ұ8#���ƪvx�z&#c����:��ǧ�&
��v��݆<o;�,�1��
ß��<u�����b6�㙭SZjS��ͩ��m�Tn�u�<q��3���;�[*�t�KD*5m���яe�1����a�������5�q�o��I����Rǲ��;��r�_G�l)1{�d7�o�2?ߗ�֛��/���02�������E�׍r��f� ���pʌ���*v��_7b�߶-�c'P^o&%�붿�g������Vcm���>/��ҟ{�������'z��Ծ��˵�ƺY��$�)�{.>.qY<|@#�t�7��N��Ob���N+V"�@�4���&����!Ikn�6s���x��q���e�(��6����Gc*���@����4���#����q��ۮ�.��Dr[�|~���tS��R�~?�,C�A�5/�(il|X�tTP~մG�v�d0���h���jZ۫�%"���`�b��2���9%Mv�Y�� ��i����D��Ze[1���*E��r��yV��AŠ.$��m���2��P��J���#���=*6���}3'��ގ��4�Ǻ��-y'{�H�\���}���@|s�J�Ȃ�̜ܔ�1R~�.x%~}�'Z���H7����2�9[LA��P�ص�=Ř�(���x:R�kx}^��z�)��`g�YP!��!50����z�����*�Ǔ��{�=-Hda�{�-�gc�!?��K�O���v�j�/��|��_�"�PXmoȬ����+����*�/��������X�/�"12� �V��b"S����O��,3������NF6N�r���x��P��hU���N;2Z�8YҹK �Y��l�ɲdz3H\�]Y�VںOz��i���Kb([�#����n4hVT#�
=���:4�H�z�t�EJ٠m�!�r��U�Pr�p�˂?'�� =!qbi�@ �yzUz��ߪ��_��o�"�h��VKc,�����~��fs��m{$̬Z�+3r6��X�80ф̀�L�޵i�8­;倓�"�htˬ�u�*��H/j�ܿ.B7w�@�ż�w�N�����s`���v��N�&�<g=���Ϧ2��J\��B�{}s��M0�s9�����(�I�l9�y��,3��C�y8��zu���5�ZC�f���Ϭ	��2z�W��a�F#��5�CO���"�<plgR�q�;f��Q���� ]�Do���
A�8C�o��}$C� ��e���@�q;$�� �}�Wcb�	e�����H�?Dn^�<L9����`J.v�1s��]|�q������iٵ�яֈ���R��.�^�[5Y�k��7$@[��U��)��#<�¾��O���҃i������!��Q`�^K�bu�j��p�r����aui�?{�/�����;�3�f���m��=SWs�Ԭ�v��ya�У��aV��A��@��ͻj�KM۝���;��3�ﾶ%���~����'[��$<	3�8���F�{�!ǘX}��{��G��?[</�F�X��Bw����ÐM�\>g���B�UjÏ�f�t���eW�&-���] o�Ld��R�t[���8'D�|V^_�����/�6���fs�&b�+�b�_%��!J�[Uз�`X?�cȫg�� Fk �(jj)
��i�鑌����0��e���>�q`#���:A���68x��1] ;D�I%��O�>۶ʢ z!�:f㴳t����`)l�2# �3�<^���'��4�7Ԛ*�0�8�O?�n��ܼ���;�oZ�o߷�"�6�����,�����Gw����~��
I��My��.o|6�/�b����c�)G."F�(���U���k�`����tb���_߃��wjcX��{�(k��l;O��GO|���M�_�3(q�z_�D~е�`��$tr�j���F\�lxQG��k5����Wr_�##w�x��[�v^��k�7�0���������KE~kT�_ZYP,T�Y�癨a8��t-q�"]�ʔN�h�w�/M�B?�#������JW[$���se�7�����1d�=a�7�7
s���]~�[�08�)7l��^!"�hr{�ڋ�j=�l�{p�[kp���}Z{��ޅB�}����N�k����9K���$�?��/���_�Đ K��y�g?|�̆h֮��<�w����ؿ�o�hf"�'��ك���0[�K�'�J݌ Bc :_v1��@5�O�&��f]k3�6��z`YMf7���b�N~M	ݟ��|@��;q�\����R���T����T�3lM9����hN��"�\�|`t.a���!Q
�+��R�9 � �(�F�� ��ضD�j�d���g9�r�k=�I�/:��ܩ���йjk0АX�d5^�A{8M�U���?�ÎXW8;�@��J�,l�x[M�1S���0�f�<A���ǜY�Z�C�����wG2�@gVmM�a0�}�4.�A��?�����pأl�p�Bo�)1�X�d�M�t�`�,\��S�K?	_k�Ml���� ���4������]7�s���u�ǯ 8��S����}�<{y�u�y��\��=��qfw�ϟ�$�n�ADn��t���'D4��z�p���#^ƢF���t�zS�*��GP����\���j=�+�Q��v�ѹ�i�ȳ���1����Gũi���m�E�I�d)�jw\�����l������5'Cp�7~��1y��I����3ww���a�6�R]K[�^��m?����{w��Yh��߹w��iK̨~�P#s��*�`O����Q|���%�*�ҽ�r����`^?�Hi'|���A����P��\I��4����
�E���L�@ަv�����ݼm�ێk����	��h�Kk���!���ݲ���NԳ�E����zQ�7]Wx�]��������m�|6�Ta01���]�8�"W�����ٙ�!��4&'ٿ�H�J�b�����}CI�E

w�=���E�u�j�h�F�Kn�� � �1��=@��K����sS�����E��x�s�Ժ���f��Ĩ��������/��#Ѿc�9Y8z�zZ>ȫKUch���$����CZ�n�)�^��/=_(���P����4/mG\�!0�����6���G0=ŰP�Z��:�o�Ig� a��ׁY[-�Ѩ$$9x�m}�fЎ���%�߃��y����;�h��[w��J������츄! mo�j$.�(�䌉(��iB�A�@�{���S4��� �����t3�3�􁆼 �/q#�TC�
~��8����:�W�E��!��TA�4��Y��e�wG�	�_^3�Se�n�P?�t-�+8���\r�������9N�n��*�PR�4��Cha�,(��U�ae��>j:_  ��ÿ-���Imq�
af$�����������������n��&3q��� �����mc��?��z�8�`�u���P+~�H��v�'������f*�����!<m���T��=�:R�I�SV]b�D�r��̾�rX3{a7@n��8*;QI=����	��ZўI������D��v�!�/�����cj^�WD��܈,QW�J(o`�+�_U>i��;�U0'�� !���-9\ !��m��D�q0���pY��zJ14ⷽ|Xhw9C�i����N�����07:/��`�F�jS*r>+�d�sւ�r5M:Z ��cZw#�"^��'������ ��ߜ^��|���T�Ρ�[H�g�[�Z ��d,�4XĴs�&��#%�%7������|o36�����_Qך`�g�{C��!�z�qto'*)����]��l��&C�&�-x�(�O���V�7hy
��������9�c�u־��v>JwVɟ�@uV�= �Q/��Cq�>+�DNE���L��os
�=F$&��Q)>-c��r�%I��{R��+��!��M>�u��w{@l�|�9s����Vͱ�����l��pcB�AWh���f"k]����x	�13ł��6��C<9\�A��>6��j!%FU8=7+�&�mL� ȃ�����F~����@�+�k�2Ӂ��O4�TڎR�^����[���'G3��k���1S���B�M�T+�6���uu��w�;��YX|����L3�)Z�{������ۅa�����78+��x��}:�L|��]~�6�%��r~!6pm��,
Ȑ ��x~l�ۂ���u�H���}��G�,I��\�5�:���!A/m2xt��Ӎ
�6T�Ԛ��`��!~(��C�{�t�|�RKeս$�_����5�7�Z�T���Ŋ
�&�I��������+�P��`f,�5��	ΰG�Љ����H��R1�����Mr�y�'WZDۻl�����TA�� R�b��j�L��q�V�j#��Xv��&��\bL�fm�N����l��N=�j���ӌk�
:i��j�C氚%v �8��N���D�G�`*L���,j#�ڧ,�tU��V�@���Y�����8��۪>y~a�81��ܤ�K�L�(�1"V�����k��o�0n�L�J���{RU�H��(S�f)�mﯙ����z�{a+�"��ܒ��=���!9�n����a�����[\p��Pw���&>ɩ����h�E,�y(����4�=k��4P@��R]?����d���ൾG�ꚚϾ7��v�`�?E5�H��?�/�;-^[���d9��9!�m�û��h,�ȝF�iG��m�L�p!�l�~��J�W��p
�� ��g8�L�b4(F� �@[m���ѻG
�DG��r�yq̟&�y�*R���l��'�+V�Ri;1�/�2|"~BGcDh������dA6lt�w�|?䮞���99
 ��?�:r��}�bp�{���5i!u��UO�ָgv��',q2M[��]wz�BB�Џc-b+�r@*~���M<r&)i���@�v��OS 1mܮ�r��ގ�@qX�Ux��t�FB>��(uIx��A�[�=ӼW�P��@���"�S���|���� S*/"���%W�t~�2�|;¼2��)
�ӊ2��S�� ��&����B7��ż/H��7��'j	'` �h��������}q�����=�Y��1�'�iß.-�.;�����<ܰE-��R�M±1f�$�4��v[�ͅn��˲��4�@�&tr�C�}��t'��m���IR�v�)���<���8����h�����OH��nYWC�)D
b�I��������|D�2(����c�ۆ�����膾_{@Y��f���}O�@�b���G)=�����s� �R[�§zQ�άq���J�+�xw�M��p(�Z3��O/ƹ�J�`�"dF耲������K9P��{dVO��$O���ۖ��y"b�S��� ^�[�`z`9M���43�n��V�u�6��|����gz�����]�g�6����;?r�Ck	MR�2��b�'�ڑ����V���f�d��ɰ��݃��������MPM�Vb�0����BZ�<��<o7�?�x�з�=��ȼd#]��nR���V�=���r��/R~��Y%����X��_���%!�kT�]�E�L��"л�7:l;�
�N�Σ��|��=�݌��o��<��8����<1y3e��9Q�{�?��蔥����x�
�����J�R��ޠ'�5�f#�=����
�`o8��FP9�LO���$ݯ.UA��z�����k?��f��Ed�l���P\�.Z��w�T���_	���[��ܮ"N��{W���KK���_��\�a�<�J���Z�๮^�'��(XE�~|(~�A��I<����(��K����������x�E���J�#��6�@F�{8�i��dRE�Dr�P�Ħ�-v� �*>���N���t5�`�w��-��4�����=�ǭe�<snJw3wް.��Z���)���0��mAGPԏ��h�& ���/r/���ӵ2�'J��v�=�[�OeO��K
܇̹W1Z�ȼ�ME������A�79d(ݐ"Ź̓���)���ڢ�3�N	�5㓓_��ug�K@x?�����+�[>Rӎ��g��f�l��e����	�p^]�G�O������&Ƶ��c��Qu�C����Z�h� +^�)Y+�P$�.!��#$���^��⯁vw�2��E�LU�v��'����L|[�w��� =us���C��t�I�8Q��2f������%��o���=�u�1;pW�����6�74^<����S������Q}�~��٣��;6�[D�<	DB��)�5����~�X�4����o/
�&�o�Z�a����w��~��~w�� ����s�'�s)�P�΃�ū�洌�/z$)�ȘZ�tV�̰e�䴠*��Z���M6�:��B��_{		�|1t*�7 �VI�E�+hS}@c�KaxR2R�0�w���,�=
5�\t��,��]����~����E�>G�'E��vj�u/~;uo��e�D���ɰ������<� wW3ۯZ��Me�����p�ގIV�� Ǻ��G���D�Z�AY@��ꛜ
q&/��Y����ɞ/B�n����q���
$�vQ_������<���+�!�����m#��/�+�~J��)����)8�h�]�����	n�)������(NO%�gV�_��@�`S�9�殐8�l�J'���$��C��+��Ȥ�����"��l�b�����5Y}��z�８�3�%(�^�R���a� ��>;D������_���Z��
d�Sn��M�V�m��ƃ��j�Ҭ[ Nuj���C�?�m�r 4%��%c(��ړ��脶�ӥ+)�-����]Q��n<�����<Ʈ5Y���+��0�Y��m�N"��U���^F�~�8%�l����b1�DN�AF��#&8�yᆺ�~2�8?f�-��U���ΊB��w�v���;-�� ��Id�@�,�,"�����&�Yb�>0���,��F�:�E�h�e��cR�v�^9+:��h9�Y4:L�����"%�dي��҅��E��q(�<v�j0·R�Z�Å&h{� H�3�!�y�%{n)k��7&�N}l��X�b/�VYçCFQ��C��Vϻ�Q��$�n[��Xں�r�͐�k�ep	�ӄ�ȹa}��v��_b�n���/���c�Dr_�u�	�u6TT�Lh�錜��3[��B+	C��؝��n��-�B��.A�wwww�� AwwM�$Hp'xn�%�C������g�{��ZߘU5gq�A����y�Z^f����ҧ��?��_�/�I{M�}�������[�=�H�svl5H;ꗶ,����ĖjG�jU^6*�\S���3/�i��m���d�K"��7�i�z�?7�~ADb�b\��xz[�xٵ��˗q�� 8��_̊y%��Z~�� ����:0����I/\����<T��(\l���J�>�dΨ#�W��$���=F��s���d���EG��gdӀ��ӹ�7'9m����)��Nن�}�p	6��yajs�m�a�Ɂk�";Čj����8�	�x<�>J����m9Tga�_����|u;c�Pbä��'��h#��Z<cӯ�ϳ��+�-��@&��竭D:˥�R?����ܰ�u�2��׎:�DW ��A�ty*G�-\]�%+|~쒢��8�Y��I�?VJ/̼��3����Oeɲx��ۏ��l��w���9��y[�)�?/E�1�]���T�!�w����#�}���5�Y�.m;����B*�����#��&��
~U�Hkq�<�y��;vm�����$w�)k)�ѥ��	$���{'�c�:���f�x%���������_��Z��S���E�Y�JT�_G'��{(�Gq���"**[Y�I?|>�A�"4����_q٭�m�����u�[�K�ݵl�������D��R�2��g���F�c3kg�K[�ȕ�
�%���}�)Ьp�ƵQ����v�~����Q�Pp��Kw���f�X;�a���;p��ߩ}����ƚ��3��TYߵMk�H�S<𔣣��FՍvf)O���}fۘ=}�H�����uԶ��t�c���_;x��:��I�Ҵ�^���e�hW�"�z�:)&�#�=9'�6��J3r�9C������3������WH�HЯ�2J���ܸ����F˹S�X6�<���N����C`�s���ƆV5���k�'D{K���G�۶�@�iO���hG��Ȇ�0�Z�S;��40$`�紴C����%�JZFf��Κ��>�����)s���%J��ٞ��p�<�R���n���d�826<
�扬fʒ�	T��c�� �Ѻ	��﹟�������"I���ո��x�]��1��L���s�luZ�GYl�I��,7�+@?/�ò�d�K��R˕J���O�[���
y����T�������hU��8�XԈ��>��6<��(��y��G�=���5&% �v���X�?6ϸ�ؒa�����0�h�|������Lq�՞��G>�;K	��U��Rsu-U�eF�Y�N� �"@R�t	��	�� b@E��M�x��'�Z��e�\ٲ�\X����k6-���9��E�T��߱Q��A}QL���9ǹAT������]�#G�r��������b�3�U��r%O���������l6�g�!�i�W��S�,��Bc�a��x����8	�)��t�s�F�F_:� �%��:��V$(~�@�"�ې�Yĵ��u�q`�Q#�$�X����QX2ǯrȄ��}n	/�}��}va�Bۉ�#��� �ptz��1��7M����z�0j7ȁ��������꜍3�رv�d�v��&	�i���s� YK^ц����'/rMt��P��Kk�Z�X:r�����-��V��_����R���!a]���JiXJJA�7�65 =�XU�-KAQ��	�6�6.C(��I"_�6g<�RN)�}�<L-�k��e֖[MMi�ׄ�~��aȹ��hj��Ǧ�"�q�<S��������V����U�����{L9�*6h�	�-�H$���>�Sl�w�7UY����5��#�\|��,�T���Ez����$��BMp�c�#�e�j\���8����ʚ�K��!��Tﭔ(������w�yd���m��@	i� ]`��[��R��j �8�_ �q*�U[c��#f2p���k�-�MހkL0�ke�	���e<e :G�z�ǉ8ꢯ:i",-�DGb�d㙔]#�>��Y�V�M�/ZY��IJ���z�_���1�#��s{���e�A
�������E։Z�<�F��q�]�]��s NT�ш��n����R}��J�1��é������kğ�E��
�n�m��y�o����f�l���c~qn��0���t�0�aS�8iЭ�;ڱa�ld�N�Ysޟ"p��A��էe3�H�'�Li'{JQO��zMp���Zw12���a|޻[u�G�S����;K��߫��
ă���_�Pʹї�ڴ�L4����9�/��S`CqA�>���\M����d7V&:ٵ�3h}�l�!���X�`θ����P۰F.��q�w��M�!w��Jk(��#��oCO����IeA��m4V�W�VA_����4(h����M���^b��6��<� �?���c��K�	OD��m���^A���?����Z���P��x)��)t�1d'BDY�?�K	���ʖ8P�Y����	B�\�;)���V�+c��2F��r0�[c�����m�09�e�D�*G���[˥�m�9e�����}�p�H��Ja��j�t��Ie���F)є�"�?�b<�<�J����\��ҷғ�_�m�bsn��Mǈ�U���"�;p�j�._��'t�sf)'V�ܣ�;+5\�I�)�HyyV���QX.LM��1^C<�y*�1�4f���s����5�A&���c���VC��ɶ���sMU�65�������V�����hi\�#[[��K��߉�í(-O-''H���q��~u$�Q����*�(L�?9m5������Ϸ��eVs�c�ͰH"���n��SAÙ���|�@}�dPc�(֦��TʬɌָ�i�q�ӗ�i.��UX=�,��/ڜ����zͤeb.-�I�Y���Y�G��<L�E�=S4�G -6�q���"�M>�lMF��W�u&��F�X2WlN=^}�����q�Di$�,��f��\��Ueg]R�	��ZGx�$�`, H�Z�\�`T;�~��	}iO��N���Yl��l��fVa�%���¹ �m��e�N�|#~��ceQ�z�z��j�A���e���mJHyа�j���m4�:������Wj�9�.��~6կ�r�EQ#�6�/����R�r�6�{�#��܉�h��\նl�_�4>$a�u�(���$�8Դ'k��s�K�]������p�qK-z�5�I�q��^�6{�⤠.��h70������f�AE ��
&����:aҨY�_�R��De�:��U�{��3T��0!�J����&g�??�A��V��	�5�כ��7���>L��|_�%N-���� nH!1�$��론�C���]�v��k�jOf8�����:�x�e9,��v9��t��xkc���ʝIf�C��hW�`I�1��x��L�P��qΐ������`t���Q��,UR�k�t��=Ӻr�vPH��X��ⷑ��9znp̣,�or�g� ��~�U*��ٛ{th9�����2z#�壹J��2�������5�`�l��8�g���%
"���0,~ɻ�8ǝ��� ����f7�Jx�
��5)h2cZ�é0�9�^�����Zƈ���@w�3�I(@=����>����@�v�[7U��F?�����%t㵡z��������ݝ�����?��Q�0��:��D��i�����9Zl�^�@0��d�n���$���R��9��붳�W�.���m��,�9�k��������2�9�]j�J�S8���A�����D�%����ddh�qm�lN<�z��f\RôZ�T�y�������y����Ƭ_C�|cS��7%����.G��Z$�꒗�p#��UUӠ ���댩'Y�Mh�P�t��JuȌz4x� �	o3MS$�u������si�����\��؏��8���]h'�<�>[�J��a����Re�@�Y9W�џ���? PN3S�u�|�V��.7��IW`��T-�5�e��	�u��#��w�6�|�� k������4D��e�!}�\3�Z��'�gv����)9�L''��#���������5ɍb���Đ����{r�#������\��H����]Z�:v���`�`�I��7�RH�L�lN���������dH�S�{k1x�3�m��/�i�.�
\���a<"f�i�m۠a�`���34��Z<�n��Z��{����H�y{��_G��meEe�]�K�Uέ5�0(��˧,��'�5s��r𒚲����/d��o��N��=[�w�¥���^3��,J89a����*��p��ܹ���x�h��n@������;BQ�q>���K�GԬ��{���X�\����~���a6�I��\��?��#O����D\�'O���eVCWD!�M�#�~��?�k0��[�@bX�v+�����9��2��y]��Y��]9>a��7�;�n$����[.�o������b�7a�n��'S��CfҐ��<����Ut�f�F2��ylR3�ǲ��y{� �sI�%]��������n c���[Ur鷅7��E�'"N$�`�}��u��&,�m#c���,���H{��p4;�)u��p$�e/ˑ��G��N��EQ���0��܎d{���hEip���}�R�!hZ�/��@B�uC'Uߒ�v�r0�$ӥ��7��[el��FS'V.0��z(G����,��wY��~�p{���@P[��V��	�����Ƒk{��u��G(T2�<���`ij�4?v�����!G�d�IE�>C�R��WE�i�o��-9I���z��:̐_s�p� ��"��}�_�_v�l�b�M[�T@�S�~���?U�Aj>%H�&ׁЦ�ColX�C���߰�|��Q���XӼ�UZLU��k��������?��KQ�$#a*��%�
};`."������uS���f?���`�0��hٱI�i���9�B�q[)��xg�E��U����$��Z* �����"X}���9�bi�7*4z���6����R��H�7fNN�|aS�]i�\��Ӯ������t�6Х�����I���ز�v��/��{�T���Ix�#�@���A����6���Ģ/EUqu�*3���L�P�Q��/�L��S��$L긣-����^r穣ks�-S�/���Px��W��$�Q�P�R�n�F�e���)-�����KI���E�Â�1�<<��>�E4�$Gxv~~戁JK+D��e��(��:���}���&�@�ő���e��h����6��`�XdÊ������H/NI,OX�:<�b��H���Ēp\!��P೷T��⍹���	��|De�.�.s�$�B�E9�Hc�Qw"U'�p�Ĺ𦫠5n��y�
��ge����dBl��1�z=�;yi��6Lӎ����$�R�<2a���a߈�qH�G{�D	ύC`�Gc�km[~s5Q,2���6��.�P	d�S]u
��U"Tɰɬy��;!^�ʋ��"�aӯ�E��nzU�?�J�<����}�օ}�ao�#|H�w��Q��H{l l��K�,V�CS�t�}��D����^N�ō��
�er5��ZbR��Ektm�{�4�A���R6��Qm�(�0��	��M��?P���b���8�-w�9�i��!�ʕT�{�6�a���5�e �8�~�(�,/�I[���Qn�Eb=����c�T�^�*3c֪�&���Hy�D4$G��&�+tWKY��v%��:�I�v~-�5w��q/���_B��#������L���D�&l�����,�u+[�q�Qjb�r�𳥵�1h�]%��:-W���.�of.l��Q\���N�_�X>��̦	W�g�A'� �@5���'�9���9=�~�p��p��?��Z���<I�ْ13��|0�[Zյ����,�i翬$yN�7�� �Y�	�����C�?0i�����,^���,X�t�|�l��s� �ݩ��"�h<�.��$�n*9E�J�6����*CЁY]�{v�rs�r�3}Y=#��N�I�H���q�5DD7�~��*Y���mkT�Z@��@�r�{��3Y��&s�xm6ھ���D����̇R<|1&j���K_�qQ��	zi5HW,'������w��y��O}]lXY�2w;�$�;F_�[���+��?n�������E��F\�G���\�Y�D�����߳���;�Tc�����i��z���>O��21��N���Qxz�%v���=g�f�M��$��^:�bI�d1�	�ÌFu��On�R �I���d�(�\Y�T/��H�S�{��}�.��Q�6~dil&�\�yg,m�~�K\wAI�,kY�tV����W8Dڦ��CY�}�3'P��4�XuΈ�xP��#��G��7ݫ�Ct׹n�����������R�[u���o��rf�ol���G�#�����H7jEPY�W|8���*K4�N
i7�:!��(�s\UuɩV�j�}��9Q��tS�iN�3�11���㕺��Y7��ó�V��\�i�X��6�`ja������[	ЙU��<�+A��x��`���𭋶4��w���b���"{��� �~��;��RUk��j�D���)u��2�sWQ=TL 3U��;,%�h�2��Tl|㣳G|F���L�=�&��Ř��0h�G���Qr��1�|������ؕ���o?;b,U��8��MAo��;�^�O�F8�,��Sxi���m��]�_z<�^��8:	���o�X�-�ﭞ�`��m�2F�O��a_A����O���B�-/z{9�m0��:�4�f/=��ԐX�ʼ������}� u�(L���n�-���U��s44<���ASqp�dH-�L8�8cy��'>x�	�Hu��v�6��|�nL��nl�S�� ��r��D=Y���E�����@�?Od�/A�� ��E�`:�_O��U����@f�W#�����:��ǖ+��U�*��������O��3 ߕpRFpN*�,��a��CZ��Í�	`�ӥ��[Y{��N@��(~5��;U��6���G�@�a|�6�f��3"04�F�g�cҊF)ͪ�@�*�P��ЬQjf��MB����\jC��QaD���8�pԄ����^�5ɴL0izd�P�A��f��D@��z?����F��]E�#���=_s_'h�$Q	T��g磿Bvps���?$��^4�0�T��N �������A�N�:[$)�ˢLcS{̿Y1���
z�o�@���?h��uRS�EkWj��bo:�L$L��Ke�P9��3>Tn���%���#�m��0^�q�ٳ*5)�+���1k0���N�I�I%B�/w�q�p�>�#u��r�5���̃qZ����Tl�k�{�j�K�tctc3zb�K�+%G�s��j����.�b�.?v���s�ǣ�����J����(E���V�
������ĵ��<w�X�s���<]��{�Nw����"�m��� a6/�4'���b�7�D0D4� �#H���$�q����ʧ�T������/$���E멝�tPs�s:�U:�ݙ{���l�4]=��(�����*%A���Ӭ�h���j��MX#��h`���"���z�E��~�տ>�������/���p@�4d���u'�J+[��B�_H5s�4La`�f�	�f�jNu�d�8���d)�~��9��?Ɔa���
���x�<�#��_�>ee��R�m��ձN�M�7���F��/��I/�������&b"Gr1�@�ݢޥ���'S֗g�}<�Z;з�%����9�d�nA��e����2 �$�p�9�^G��x�ep�����e�ƞh��;�bL���/g�E8l��j��Yt��[�hg��q�����-���'Q�V���h��#k�G*;q�ٸ L2�[:bJ(���v�1I5���Eک(�K �$(��I*4'��H�6f:�5T����\�m��-P?D����Tu7F��9�~����v��BS�q�o�IS��z�5��?�|�}K��vn�+��1�fM4�?��Z�K*�����C�VEqH�C��~����,���y\��G�����Ȳ��0�#!maf�s��qU:q5;�`5q�YW���-���&����E����g�,֗�̄.dr��n�h�c��m��8Ž����ip['~=�G��֠���h7S���cp<>ut]K�X���g�C����X��Bչ�FU�~ֈl����7�.i�x��<���,A��I�;ɑ�'��6pU'�Эp �;�j�sۼt��`1��3_}���|Rhh9�WM�ɢ�q+��>K��"�R	� i�v�>���O��&P͞=��1�%��*��]ٵ`u�E&h�y��ID���%�32���=�a|ys�j�������y< �.  ��}�X�h�d�2@*~��0��Q���"�.G����}�(V1v�qЄ����y�� X����Yc^���f|�Ikj�[�D0��ҰN���Ev��Jշ�d`����ڻN�L�Pe�v��%ϳ7M#w0OJ!�4[�m�OS�,S�[�s�/_�����V΢,�uP
��Oc��>i�T=;, ��z<$��z���a�#C�xR��[NV���7[��_���gm����^�,�O�Ͳ�W�<��Ȋ~��NO1��=�dg޴��>Փ��d�{1�$��f�j��ڣT�������GC�TLCF�_$$a��-�����fu����1z��~�8Z���!K�+��x;w:�$q-5lܭ�8d����:��FSd��9&w��Hv�^���\���'/��\�?J�ٸ�{s�c>�o��~Sv�B&�� Ia1�w��@����	_!���y_�V���&�#�v6p�Q����љ��g,Z`.�cY\�fda��Չ<4-]���'��AG�;�i�����=�����،�9q�%n�O��c}ߧ��t�n�z[���eIP�J�$F��=-OتUf<�.�K!�}_����⚱�?�S,�z<�>5���7r��Ij��h��D�&j-�G��&I�]�Tr��Iy}k����T�[`�T�(����xR�o��d�~1x�6����@Q�� �f�G�?���r�Ma���J���\f�ۖd*�Rx=�k��ۆ��`�X6�s��d�b��qC]��Q�[�Ka���0���<��F��0$��6�?=@���ɒ���z">ZظZL~f�fc���Jh����R#=ehH~���r7B�{��m�^�ɧ��700=*<M�����!��m�[h�OlQϣ��(`&`�v֎S�f�o�s!�(�-¸5ʌ�hzAa��,��X;܍
���z�D,F���'���oUmx�?����59���6�09h�����R>���	p��D�T��m5/`�N����f.Y�k�J����>dS㞧��r��Ț�3L�4�q�br��`�%υ���B���/\m�w��-�~�s��8}������E�9��~��Y�|�o�����;:E��P�J������7�?�~���q��iox����}+�����	�ND�T��씜L%B�	|�J-&J��M]����g�*o��D�@\��tF��c��=݆&xݦ}�z�%�T�k��&*��^u/�g�#TP�W}���U��Q�C��r'�	FWj���.�M�$����q�C��[gB,��Z�}���U������ah%��+���E�Q'M�^�ml�[/����}�'�=�����0���H�P�.��3B�E?)��S��n.�V+��b?�7��O�	j�� �d:Ō,��.̷�V��p�3��G�ņ�#*���%7wb��T���&��|�H�^�j�
��\�(Y-�ԭ,��pe��1KFx�M{^��^�q�3yI�,�?�2���!F�{%� k�/�좶/�&����Lȍ���a�(�%nǧ�i.7��g���<�I�}�L�S^֭ZA�G,V��EN����p���E�6��4ݒI��8��Ω�E�ԯ��?W�U�R�6\Y�Lg�Y^�$���|�C�����V�� ��k��J��T�^����	2E��a�K6Tg�?�T/����� ��{�2�,;�e3�Hϻ����&�'�0��Ǎ���y��U�F�6j��X�����u�6���b�d���N�-�&��58,�ѣDqe�2�N�P��V{�dN.S�	$����K��tcp��N��f��@�8��@�o��p�}}U6�������2��̬����p����Qwo���V�kA�?}���a�2��L{�*�k�P�kM���YfQ�����䤲�x����kϫ+��P���d�!�*>.�����
Zw���A{ρ�F�[� Շ%Ii�kėN���t�*;�'�|�?�l�3c�l��h�����`�0�/�nQ���SuWC���P̀N��5PG�P8 3�U!��8^N$��a���	����qǳw��F��]�
�{oUee���}>/4��A�V,�:�QA|S�N���t�w�Ll~G��a�uU��'@���D������^V�T�����n[�8�w0OOM�Yy ��g!f����ȍ?�YvyB��mVH0��p�u�]��O�UI޽	�mـ^�i�8�U��O��1���ŭ%��i��=k�;u�J9^(�>a��Vޢ���/�&Uk�<����T���Έ�b�y�x	1a�G:KoG�-�L2P��|@*�w�IA�E�$W�P�'�u
��Uq�{Z���ڤ�FT��b�ِ�o�_�;��&8��t�_vŏ5���F�Z��������>���o��&���y��{�PM�yXh�ּ�|�b(�=C�K�ϴ�8�N���2-тF�����tW�jhl�v�Z5
�RP�����;O����z<8!����屷�����|{zh��1��������a;�O�D�E���5��@�キ����/^�"q
-��Y�an���aB]n� �7���~ݨ��;�S�_���8��3�Kj!-�:�A8��Hq��	}w�eS½�e	��'|.�Ý��b[,�D�<���|�𯈨
9Ďs壥�e��~F��블W����� Ұ}8V�Kǻ �T��]�~5V�|�{t�ذ�D����(w��j�J���h�ͨ<��lf:\|�x��(������xG��F�wM�Mh�~�1R%�r��E����H��f)|�����SWuX��&9���}Q�������?�����+����[mF}9�U�Ȱ�*<���(>����~m@�dm��Y�	�#j3E�4z�dh4&_b�$�]u�\S�7�&��Wm3̓��r�`�n��������&�>�Fk��ڕ�Yb�ƍ&��al������H�?��nOKs'� ]ْ��DY��QD�v��.X�8�xJ[&�������P�����#�e�S���h*�Ck1j&!�7�12J�M���L0Ye ������o���q�e�s%q�\�}�v����9�/�Mݔ��i}����(�<v�3�Ѿ�]��-.�l��2dn$u��SE`�8$	HƳ�p=����	> �zi�iP�Z�d@�w��1z�ջ��Υ{,��-�B��wj\(����6���q� �J�c~���L�oM��a�%�gf���w���!TD���χ N�'(��9nņ3'L�(�F�)��[c���<|cݙ.E�?"ӭa^�z�=��i`h�@�M��H�~�� ~�ƛ,w�ý̙D,�����z��?���l�!�VA��צ�Oò]�s���$�������I�;�I$u�P?	@U\��L�>NL �^bR�=���xk?��T����?�3�!�N�/��w���������%����,6��������e6`�5�uq��e%���䔕�Z���d���n�b�ϖK,c����]��j?�֡P�*m�p���&�<�H(�}u�	��ҌW�k�z�	�}�_�X���#(�a>��]���*���\�9^WT������^�����K}�G|���S|����?�=�����4��Y_p��YS'�����f#^rRIw(�/K8_ ����JX��{�LqU�E�n�U��F�o�؏ ؁�8j@�k�l�P�0d!���I���.��~T�̗�h�/؝�� �Am����7�ٚxN�?�7d�V?�4);�:ʇ�9k����S8+��8�������ZY��Dw��+F$���۷ـLL#OƂ�Z6�;v#���y2z�/]�%���?`,�^��ʢU{e���Q(Q}F��a�f�q��� �x�&�*��l�'��6Vr��J<��[�)�/��1E�П;/����UIi���L<��ڈM�GH�nn�&�ڑΞ�t"p��n�-�����Z�~�����3]�*�æg����%��L�C~�=��~���V���I��Z�+�3����ˢD�k8�ln&�6����/������Bմ~�3�U�9�����e��{�G5��g鷗SU�g�pfm�FБb��1r�!��b��Ȟ�WR��	�
�!b���D�v��ٿ�Z�)�_���&�"�bBS>�Pa�\hs3�s��V�b%��j6��mi�E5!E ��]W��i�(ûPڐ�~>pzmX�r`c/��p�kgj�y�s����5	1��ӱ����(�	u4�2�R���bv����L:ȥ�h�E�
�au��eM�΋���U�.�׀ȡ��Ss�oy�#�	�/�^��+劙�'
�}t��qH-��/;��p&��J}��2�K��O�AC���ʷ������),��cD�<d939!�Ɠ��p�J�mRPy*�x�	�Mr����N˕��:z�݁`;�Ҹza�s�1����䐌f�S�U��O�t~�A�����~���SwÏ��v�$�H�?�u��7N��o���*�rr�P���)F��xYX1���� #�+}��=O�A��������~�0����|��9r ���BH�1�����=�'�Ǝ@Y��a�xR�;l���@�m� }+�T��O@�U몚T�F�.�Ƈ��f�Z����n�f8��Fz�6A� �h�$�Wj)��{�h+�k�H�*��Y#�7h����ZX*�	+/�-���w껻��Ă�����BH���<l���u��V���i��b��P26��EVq����)����k��)�X�OCd�K��g��UO��bsqr�ӭk8��0��͉ށ��x)�����Z�K�׬1'*�������v�dkS��������9[�榟�w�9hP���w��8\�w���B�T�L�W�����[�ѭ�V�s���O	�:�Ք�N�}�e��d���,q��d�s��:r`�g��P+�W�%���
h��1sTT?\<iNi�
d;j۬^�")l���QWx��#��C/�Υ;C���ě�
*��������]�����`� ��y>��*\�m�0�d�r�����e=D-�H�nέ���aSjE��>���fB�YZ:�KWuz��Hc��3�Tk:�ŴygQJ˗O�8C�^�φS�̏�tc�PI���򨮚ԑ��M"d�7B�r�S@/�.�lkG�	k��f7|L��,k���^�Ws#���i�j���[�Y֙���wBz�!��!v/$��`�����r0�a3f��,���*RՄ����xv������tCQ)�uIFKR4$���p���{:�b�+�n's��ѵۍ�b�y5b��Y��Z[�j�G����[��>�0���\3=������>|iMa��#Hc.����h,Z�����w���z� 8�*���̫�ӢK��̌��Q�l�>C*Y�������y�ɣ�B~ �e۵����R�c�� }^ԋf}�ԕZB�75i5s��A�ujH��~>\�feJ�����R��d�q~;�:�K�t��y���� *Բ<yO���+$G_�v6m���0c��ހ��~� ������\�b�a|�G�;"�|]Ĳ�'im^��!X���#O�Zlq=�~MH��˥fu~�2"���;L{��d�5D��⾨7`w�u��!G2U�����9��%���&d�]EA_F�vE,�"d�D}eFuq�۶ɘ�f&䫾�u,j���v��|�m��V���
9t1�(㇊$�`�|�PU�(9�K�Χ(|L�k]�H �C	�MD�Z�t���:��B�ު��A߈~�t���������GOQ���z1o�ArO�,�B��u}�6S<��g�D:|>ܾ\���H��V9�^�a���A��-1��7��xQ��u�d� n��2ĵ�A��rܓ�2����fT/�j�]˛����z.�<��l�&l�2NG��Z=���f��0��v�����*��g�)�G[=�����Dʠ*��I�
q,���8�g�WQ���Uh��XH�BS����%�Ѩ�*ͤ�{۫�(i,�s_A��%�>l�2�������J���4ʖ�ͅr����7֖�1Bf�(j�N�`)"a�Qw�������_T+��7�\�emdEװ�Uj+)J7>�>J�!���K� {�Z_�>#��JB�}�F5���5p�T�J,I���ԧK]�l��T�%�%��c����f��S�tZ\�}�V_�ZM���y��<�`�W!g%�0��Q:��o�e:�~x���dS��[-M��ef�9�oQ��Y�S��>��So�/�*����%�C��i��u�q��%/����l����@k�8e��ʝ��m�[\����!G>JAx�������kp��3�!]�[x=���r�a�XT`Hإj�7�x(_|%~���~������[���#�$J�[��t������c�%B.���g��c��#tA�W妾���2]��i+FN��8����+�8����cm����)�?����)|C�:馃JgG�Hb�L��f�WT���� ���=��$'�e�=�L�)��P�O��� ��"�����V�?��	~����a4�焸%���p,�)�_wpv���ӵ5�NhH�`;�[����w�Oz.�/i���֯��,�(������`$��s�YM��Uȧ_�k-� �<��T|��}De@U$�M��h1�P�{��wU{�0�f��o�QP�^��<$����J�ٌ��h�{G�ߕ.��(\����Kf.��w0��yIɷ��0i뼦�=�87�@S�'�]M����O�S�iS�N1bLڷyA��ݱ#�(�EЙD�ys���&�xU!ym��?� z��!f�y����eIJ
w�FM&�f�]HÍ���+���B2�c�$+]	.R8S�c���rN̯�"�Y��!jZC�0��=0�?5Sn��,��H*�1T�u�h�D_���e��BpMK�~u���a)���N��JY��G��;jc�y�y�Q�V��y��>:�V>_>J�δu�����Z�
)��~�7�Z�2W4F���wmV��?� =�Z�.$K;Z��wP;N����۩�lO�����dC1�=�:縉#rA���h�9�A��R���fI#'�9�������9,�Z���!a�&�����R�3�R63�a��֣$����Q�q�Pq@h�@�;LO��B��(���4ޘ& �!�x���۾p� �p�J�~��=(ܥ��L� �!I�"qLm` d��{�c�Bq0O�v�0C<�����QFUC-V$��G�7w��ON^Z��.�윶��=�F�FR`b<��0���y_ߡ�������a�!�|yl���ݳ�����S�"�bM������zZmb��4EF��Y��>U��4JC[$�%�_���7�&���B�8�{E�9�����%g���tO!<�|����7���
��%#2�	��F.��0�8��q�$U[;�ո��e��R�!�GGڪpEn���-���䚦�T�Z��
�F�$K�����i��p��s���Hz�$�=���5ˉ>�OFVm���O��p��j���e�RD_�}'����_�����̮ݝ�U�$�"�I.N��`��4�Z0�%��2Nm�%М2�8�_L�݅k��� s���Bo�PFBl��Y�a�����{�\E2*�Qsif�!&�b���;r����A�G�$Ӱ|����&�
���H�_�_,��0�ѕ0Ѷh���QǶm۶m�N�v:��Q�ޱm[����=w�w�ׯ��&�V��~kȇ��,�H��=�wgG��"T�c3&c.�:嶡�`��m�l[�x�d�0:�t$p:�e4�� ����`}>�.1U����eW����Wn�t��ga9*]��gB������к:jC���oa����ʉ�@=.hE����_z\d-�����2�]��X���5!V) �V�6>�;H�q��_+X�x�odlu?diW;LqklG�$�m��>q���#%�g&3�9����;E��xYc`k�J��eG�k�w�-���)����]I-�Q=��Lbj(W�e��:Z3��G��<��%�E�,f�Ƣ�;<t��%��O�3%ş�dc}���??`�T>�Xf(��)��Z��1=��C@b�XL�|��r�,�$�ѷ���͹�Q���z&�H��nqQ:�*��G^����}o��S~Y�W���c���AĆA;ܰuǗ�_8��%{�Q�G7j����u�0x�V.=8:������ʬq�#)X6<��s��3���q�y{^���m�k,��Q�&�(e�mᭈy>ޘ�B,�L����G뾚�&VV{�Fh������)v�+�-v�Dw�O�E0Qt��r!l'HCjj�����Ot9K���}�R���XK3yv�pP�O�@p`d�pJF��z�&��+bM�mE��w�4��"4��e�3錩Z�Ch��U@�	�,W 
Q�-��,Z������[�?������͓�o��Ȑ�X��T��SZOتӇ�s��
��|c��rp�����Fu�@W7ijU(cS��H���m5!�u�#:�li�Cv�G���JS���#����XAB�����u�`�]��	ʗb�Z��Є"��D���I=b�NH�o�Θ:���@J^'
���G;�t����d�R8a��S,@�׸~t�4L=� �@�����-�`��-��Z���	yL#��3m������i���P�z��?��5�ɤd(WH�7�;�.����_�dc�p�8��X��5�]����'���1�B�}��f�i��'�;u�{���}��b3�֒�h�w�uH �_>8���	N�,��X�䩁���0)��{ȣ�K�����&�TZ�D��}���h�r�%�:�����C������Dy���W��z�����%����J�ې]���+5J/[���J��7q���%)ZI.[B��R�����j��v˃�ڛ%�}���9Y e[�h��NO�4 U?�X���oK�3��j��Z �g�sf�,#��1tM��|Qr~�R���h����ݟʫ�����Dy\�wF�������ʄ6�Z�<��3'z��Ia�i�ٳA���vF���:Io`s�!9���ňQ�+�*���Ū]ͭ�w 5=ɔ�����ˣ�jL�p���<���Zq�N|�ܜ����o��#0�� ?����iM��E�����Y�?!3݀���v��|��` �q�y��=�S����A�dwzĊBe��we��r�('"WeJ&�D]�N�L)��@-tm��]{4^� �a[�f�_�u�s:W�8�T���v.���d�poٿ��n:0�Q3��2,��.�2��,�������`��Dt���ɴ�14��Y�%4���s�ۺWh(����|�GxQ�U�Y��,[���H��6,�����i&R�7�=�ӈ�V
�N,(�K�������Ł@���7by�%3gdTc��J������S���	��
�j֎StA-��Rz{�Ug�qXI�1+*8i�}q��K	>��W��Ϩ���'>����'`�I�$N�6h�)נy��e��Q��Ƴ�i;�'��t�#>n��M���c����>~�Z�.2�3��s��n��v0DB��'١�S���FH�ㄺӣ�d��P� Ջz$�}���	YH�+f�I>�U9E��w���$��y�h�#ɀj��r�\y�)
���
�j�1���H�)�O���Ga�����G�x#S��@�T�2Z��/'��6��MG���W
���}b������(�rs������u?o���Bdt�nr�id�IS5�q��o�:z��)Go��2�̞�T<��:��:ī>��w@%#�&M?aU䰼u�PHH3�ʕ��$����>�.S
`�q���M�.���(,�Xs '_���T U�"z�DIB[y�)��E
��2�����s�*��c]��PӚ�`�&�ep'i���Q/qg�&r��H��Q>�eq+��*D�=)S������\�2F�/�5?��1t���j�FVzn���+|P|��qMj�t�[_���\f����c�����)��4��Z�M�:d�c5��L5Kދ�C#ɺ�f��GW���T�dx9v5k�e�[J��ϥ������f�Q'����M�d%h�N�m�V�kEWf5 *�T9Y�G�*��<�\�X�hS�e:q��������9B�!N����P���ʶ�F��_�6M�d�Z���w�`��0r!(���4�X��S�ҋr3 ���ޓ/����	z�
�ݙ'P!��+rQm��:���u�ޟ��/0lsXd�n���>�_�I g_��a��ʹ^ۦ�+\�9{�c���=ĕ��~fR�٫ٚߚ�`m�=�.�&C���
j5�d-������������}��ڋe^c��<��<�5J�(�)��1⳪�7k�f����7Ir�p��� <q�e=,��1�}��C�\>1#���������F��|��Bq�+�t, �DFO
l�H��!��t�RQ���?i5 ��܇s�R��H�B��t?"�"����u��V6���e�Q<����*�0{�ϧ^c�b���N�xO�' 3^��\mP@��j4PԿjT�U-x�`ʭ�:���� 4Ry���gT�u���mIq�������Y�V��M[�E7߉�������<�8旨�[K4P� �B��X�A�,98�Ƥr|~O�H��0y����{r;�ѣtq�x^C..��&
4��0�[�݃\Ϣ�X[���My�Bj��	�0�-��V���ۉ=,�Cٟ��H�D��#s�E��)�'X���`q ���Q������)k#�l4r<���<�u�m�Ma��`i�`)��ez�����Vpg�5?��i.�i�_Κ6�5l��a�|K�:��r��˵B�gpݢ��z�Y�\��SMt@��z=�|n�I� b�*�@���	��v����Y>_�p�1���y�a@�� �	_�?Di�K&��k��,~�2=ԓ����[i� ��9�$Kb�.j�^�\#vd���S9:D�&��� *#�t�u�i]�~8�a���"�����v�������N���F+"x�R&�����V�J�Nﷵ�-�vĂ�3��P#D��
�q�o�H1�"�)?*4Y�=(�0�F=	#R��4܋e	nkk ��L�1�,������&��92�}���E�=���_���;�Y�.���|c^e:\a�KM�4kfL��M�z���5�@�P����Ӗ�*u[0�tD�:��.��W�K��(dG��( ����1@1A�"��7>fY����/��l�n��H�nY�ˀ��>D�c&a6�k��WX���$[������u=�H����>�|���Fu].A>fԁ�%����aM�7�q�6�J<���2;E�����d��ŉӗ>�'�����Q�:���Q�E);�]��AVy��&��g�-�]����� �H.�Y�DW4��HѾl�:W���0��5"A[ռ�K��Y�Jd��A�h���`�1۝	 \+&��Э&(���q��ͿK툿+�1���3��5�5%�5B��n��C������ѪӐ��E�J}�~3T��ÎT��U���9������/�Y��=u����q�Ҥ4�����ݽv�`J��c�y�a&�ˡ�����L��oy2Rކ���xV���ؑ���l��HPӆ��*�"i��P���X�
��"$��}��X�xԈ<�CGC6�G\�O��jl=y�ی�������n{n�ĺj3�O�~�H?�>���� �CE�3�e�U�6n/F�№5Т�Cc+V����?:J���-�痳�%dG��G����:��i��NBx�^X���pm�,VS�,�9�Bf�7��~���8%P RiPӼk���������m8Z��In��b'��Ĳ���RN��V��u��@]�l��D.�A_ E��h��_��C�5Qz}��#a:���G(�ia�
��5�h��,3 ��qe5P���V�$T��,~AE��K�[���ņ; ��I����R�/C�~��&�h�L��X�Y<�C�,���iy� *Pg[��;�K�ᯓ,������T�$����&y���,�?�8�{[�d����R��'�>FP��>�|�� 19D�R��N��-� S�����j׶���k�;��p��F�9T,����E��ɽBT��q�բV�(�d5ݴ-�f;��?ZG-�@p0�\�B�?([��n�0 v �#�Q�*���s��揚��@�*8/�P��kL��0V��zg�z/�Y�L�˥�g�IP���ܔ��$��p�pهwaAf��@�f�f��?����ćRG��zM\G��3	�H�:N�$�Wk�9� d��b�WsA�.���A3�t-�`R�	�������k�ܻ��8\C���q�\��5 %ɫ5�3�V�P���5r�A����ѵEp��;��M��ܳ�z�LD��\����\TIBb�@��*&�������	Qkbn��S�t}&���c�)�~�Q�uv�X��l�1��Wa@��,ݕ�Fs�V�n]�S7R��Lk1)��[��˾�;	ޣҀ=�GXl0�v���$s&�N��@x�,�л�@K�}�����:ě��WB�@a%D�ԝ٩i���w9�zYF8G	���_���@0U�𾂀`O�A��m�\`D2Q��ɝ��-�S�OG�á�ߑK;>�1+�����Pa�������G$U:�4��;��GRf
\5�=���uǴ疊��4.���V�'�'�j����n��:f�f�4iğG�)��*]���I��ڰq�vD�ki�`�}�����"�[U��*jʄw,H��dX݁���9bu1�c9��5	�����s��\S"�}B��ӑ��|o�KkvD�چM~5�{�7U������$�
����-�l�0��0;���̽;+����(=�E�}=m$�t}s*g����O���%�Jy����g��7��� ���撢m6�$�Bw�-�n��������	�%���(�ֺ����˚0ϕG�{�ۺ��|x���mE|��+��QŚM�P���faS���/3�smH[����<�7�Gǟ8��M�_�i�]�t{A�>C�[�Y�.ԫ$LV�e�,𡲦_��N���ۈ���8�D��N\�$ڡ�e:��}�0`��$��$$��Q�i��C�7�"n��l!)���k7��f�m�2��1a}?~>1���}�E=ٖl�p� ��7�H�[�����=n_�I�Tb� �-<{�	ێB����漂jY�i7�T�;����C�/^_���|.��Ϧ��F/?s�X��u�d�_7�sT�v�ZHU]u�:�ԨIN!h4ʐ�(p�����'"( ɀ��c�ݾ�=	ٶ׮��,:ܿ�|k��s�����Z�X��<��4�x��mb(����cQ�c���N������N�*�P�|��F��m�C�.Q	� \?-�╋��b	zIu"��}��\��[N�W�7�g�aBj���B'����ה�pW�;~K?�
���ҵ����t?��#k'��Ǘ0^mG�=|׮n���삢��J�E��
=�K�E���u��v�B3��C��st��CT��Gؐ2�xڸ�(/�Y����t��C17�`�t�t'pL.F�ҳ�)Y4夝��������	���T�u'39�`�c������Cm�,���GEя������y..0�j�@�Y�n�Y�~�~3�x�<�����o6� D��:󿜟u�J�S�R�v���mwѲs;�h�٩K�x��(�x}�qW����ô�4(��T��,�K�Is�d!o'�`n�.RK�}u�M}�_h1A�a�S�i���¼���T'��L�CSM%�Y���z�:ÕGm �f� |Q -m�2}�����Q,`b�um��<���q�����P�\��b�þ����P���"��I'����RG���Gg���[H�Û�!#��s��`���Dr�y�A���)�M�h�d�F�V����R"|�s��3o�UZ`:u<R��s��(�2e�I��3A,B��$0�K�Z-lr"����{��
K���)�8=���o��Z�St��o�Z&��A3�:�p����6��pRǄ��x��m� ��h�;����K�����e�`�ikZ@�{����;C�)~�:~����5֥�Â?R�>���P�2�pf���¤L�n�Ã�up����؎�����|c�|�Co�Ô��̔��P��5��g�Unuǘ���f�W��Q�e��fl4��o�`Sh$~B��=�6�5�B]T��PN��>Y�	�Cd����X��~‛kp��g������}׌?������t����G���Y�����_�oW��-����KD]��� ��S&�Q�?>P,�~�ǲZh�"�c�{����L���c�xx�97�%vKNd`wWϩ�=����5�-��n@o���XW�r�js�+�Q��k[��Ӕ��5kҹu��#D���Ȳ��Oۭ�(�X]��ӡ��q�8
O��ϔ��v��p�ux��'�	�b�b]��=!�gqo����k���q��*����$�٭�9u��ADQ��C��T*y��}C����lk�f���P'0a����nf<���[VE�3�m�G,��F���3�ʪ4K�����I�`�z [q�a6e��#)��#w�;p�Mq�*��4�he��8?Z�k��G�[�(�v���d��va}�.���Vn����(I���w��*����r)�l%�lSN�Y�*2N%K/�sN��N�2ٹ��o �b����ٔ���T�-��X�m��ť˯hS�`��ӓD;xbZ&��4m��|��
����x������Q�o�������!Z�kT�gI@#F��צuFO���m���	I��Ő��g�����w�Uj4�m-z.���6>d���A�������kH5'�Z/;5�J+G &����s�2}��m��l��f�Z;uɛ� ���!�X�: ���!(��N �(%�ou���ڇ��'���u�?�����������7u�&����YV�^ v�*�[�)|By���c�!~��.y���h��>�״d���E��g�3ʉ֪�;�T}�i���q�9�Vލ<��#���R3Ύ�s������_�t/ߺ������q��C ˷X]�K�+��\��0 �sg�j@3 ��T�T� K]�=�ں�J������&Ȫ%�� �.�����֖�	��'4**䂒~8�َ�c䗶��uS��oI%��qֵE�Bz�e�����q��Bٷ��]Y����!D��5o�6陵,�.!���C_��'��N��H��f�k�
��
�*6R5��ל�T���$�ϡq�㨦K����d*6���t�X�3�m�8]N#S��È.���2��(\ hqWl���I�Jo@6��5�k�FRȡG��b�@7 ����@H�����ޏ��_waU�]A�=��.9����Өag�e����L�ڐf�}�*K��>��������v��vz�?���B<v��T�@U��s�7��n�b�q��̝N|��b�c�EkC�z&j�6<��/���iդ6R++*߹Z[�x��ٱo��H�f��bJ.�s�M���g�!�/��@��~�ؘ!&�����~��������O/������A�j�<�_���B�ގ�S���¬�;���p5}X��`���"�}oo8C��`+і&�%2��7Dƨ��1E(�ؼb���nJ5#r����� d���C�����~*���J�sTQ�J
A��S�K@��Bi�FJFo����0F�4ڐ�34�	ʬ�Z����@_F./-�	�u%�R�C����Sx4	L��8;����:�����Y΃v�Ɩ;��n��QC�M!�s�%��.E���ۑ=f�M�1*4"�ٝ��F/�%e{T.�Hd)�ߐ�2�D�@���A�yQ�3�Rϰ�b�+��8Ay�#��N��>Lg��@���k�
N{�e�nZ�]nk1+Aٮ$�JZ1�s2��j��6���6����&[����;�ї��C����d�o�bٍ�/(���MefH�h�B��`�����Ap��w�֍�a�����K<�G����̤��CZ��m��÷�T�TH�Z��rXĸc9H����[��8_NS5.���]%fk�C�}z}�>�R�e(\|Ldǣ��3��/�@��̧�����:�M�7�4REa��_Go���������
.4�3/�t����9(����o���|���Ǔ�Ek+/���z�/�ͼހ�2�c;�2�/�c����2�^y���^�kWAQQVBB�&#77�qz��!?`�4�e����r�h��e��� �>%uU��І�V��'��q�u�(ڄ�#>��H�Jb��?[�'�&%�^��_�p�e�~3��rAX\�j�Z?�"�Lv�z��%K�
w-d��'�����w���izܮ1��U�b����>#�%V�	HJU4Kx-�	�u_�	��`<#�ְ
�^��S�E�����P��`�51"8{��h��%��Ŧ^�7�%��7�~����S�n����m�o�V��Xt4t�&-����W^6��N��Z ��K��"��,�r�~���bhUDe�������﯀!�+���䊽�O���h�x���觖�������؉��X��߇�@�� ����$zznHi�!�Ew9��(���b� '$�.�A�n+��Z-���E�:gI�����!Vr0����>��|e�m����������u%�uur�ʘ���w��~&�זc�>vYH^��u�	���c8y���(S3]����q��$'�Y�v�tK���Z�#�\|�68�r&�_������]>��W�2mj��P�����Ku��3��G$釃���7I	����5��/�:#���W�#��g�b�:��F+��M1R���%FK4��sy^VL�kM7��^��.�F�m�<�ak�Lh�_cN�W�ay\1Uqs��� 8��!� �kp�q����R��iybev��*�F'|H>�L.P���O�giċ�H�����y�&V\�o�R��!n�ʓ�r{ن����77Ž�g��?V���@-Pm7�p`XK:� ����T���D�����s�c��HH�;4��z�����z������`��=�c6=-�
V����p��� �YI[�<�o��㸤�5�Q��.9 ֶv#X�9����]��}��	:Bw���T�����B1��Br:��SU��[�
I�L�R�7,�Z�iq`��e�cz�P[.�4��i�~�7�\.eK7p0�o��q����)/�#j�:ˆJ?s�z��_�M�un���uA�t�g wKΨ$0��H��},�σ �5>U�Q��5�A��Ǣ�[�_�hE�v� �h�L�խ�E��+��^�
��ҀQb��_b�z(8�.�cE�C4����Y3b���	��@D�m���+���N�Q�XZb�Wc�վ�K.iJk }Z�n��j��Da##�Fh=K@����O���
7gk�1/$��+�c���a�)+����@�)�:m�|E�غ�g���M��旽�oر�0lh5�i{6��V��t��cU	��W&*�p����l��j@s�Qz��-�hoX�t=�X�~�K���z�$3a�u?14S���X�C�-�������Oi��w�J����5QPY�Yq�e'�~�yU�y�Z66F0�m��{����?
��'~m�?9���Fe0x��(ήk})wJ�XW�� J�_X���I���;���h���g��yY�_A��ڵ��n���Q@Yn?u�i����?�'�r#^����ܽN1H�S8������6,��",�y�;?���Q�y��U�;N�f��N�8��6V;}�+�ޟ5�m��n���3�D��SLA_��P�ft��~��QX���E�|
'�f��]'��}��(O�nH�>����V��(����?�Kޱ$��F~�H2�q�?rM�po�9���(ޔu&
��.Қo�m=���lK�����7�F�w"O�}$ch��"��5���2M9���o�7u��ge0W�,���i�J�jZu�!�J�SX~Dx�	�;0Ĺ����?�td����8�?Lc��t�`���K�� ���o�Di�w�3r�����uEl6/~���I��I�M�0�����>���N�м�ul�s���@�
ʏa�d�,�'e��x���Tzaլ����hhj�^\��P�����Dܻx@�XN B���&|�4�%�v�5�S�b���)��-�����>J�o|��<����H�cN+D���
`��\�\tKx�ۧ?�Q��;
�ſ�tM����m��-���=J�ߙI��EGY#8L���½�N>ۺ��ˠ�:�bD����$�z��%��]g:�iҜ��߀��'w��/N�]ag:��������'d�p���?�Z����L���N��W]�8�?��J����������y���U7����}z5�#R�����Ή�^���T���a���mG=�e#��u��|�\͸����y\���u>�ޞ�^��~�P�^�D�5;��0��^8��ە
u�����>P�:����;��1m�֊�������}L����V�Yn�lW/�!�沱dכ��p���m��~Q��F��p�_�=���^q��	x<��79��F������Wy�q�$���w���n�GlkE��&��f���0x=��g�DW�w��?���r�\����E�����/N�WW�}������)H)Pk�;��;�w��?׶���Ts�O�ԡ~?����z��z��Α;G��Z=��8Rl�95)g���6Z��K��/9a�"�L!Hp���JMo��W����l"%DLΘ�u��k.-`�xN$QY�R|pO����t�l-0Ho��K��'������Re��6I����M��UDkA�	�s��X�39H�{��\nk�t�j� [����1��2��_��$z��vYh��H�Cg���
�~7�X`��@MLL`�^���`����;��r�īZNG8t�<�w�/u�z�<f�
�o�d��W�?� ���$k~}�;-��5�һj������wx�2���k�q�}��n��"�"˱^�����cei\9>5¹�l��fgr��x^a��RZ�����$?Ѡ�"�9w4N�T{�L��Lb] ������S���i�uS�~a�7���e�(p��7�E���u�^~3a(l���s����T� �B�*%XA?��^,��\�# <���;�v�7�o���%����g���w|r��n�mm��c;�=���iW�V��'�;���9=�%���ɝN.w`����)�(��|2W�o�S/��oo�����n�j,Oث������������j/�z8�3#��������8-<�]�	 �2c�i��~��,�4'J�5q�Q���~r��#�ݍ��{(�Y^������=����s���ti y�Lfs���.����~ɹ�(�D �q躅��>x��<���둕QU-W������}o�V��m�
T�|6�`�������%�/<,e��TұP��Ӆ��a�a8m���>�J�+}o܆�Wpx�����Ģq�z.k�O�&��ذ�+ �+}"� 8CC2oy?��*���,Z/v���+bز�=Q)��f��]��������\�(,��/��3wν�-���U*�Hn_�����g�����O&�>/���n�D�B~�(�BPU�HSVɛ>	��?S�ŧ��nM�f��-�fa����� @���l��{s�VN��[W������q�ۅ���x��(��+�b���	1�����9C���6&���08�����7�S��Wa�c��z�4rdC��Eլ6$pfZ&�ȁS�.�W�_Sg�JI��	9�056�\N�e���],��=(O�{(\��HA�X>�ν>�|�	�i&��3{{`����T��N_23�^��<��!x��7=��'�ˌ�Z���f;��ƮCZ�����J>��*��	��o��%������)�~:J�}Bd����$-T�1v����z�f�iF2n�]- ��Q|��1�S�w�bPִ��!��oAD��$��▌��eq؏�$��ܒ�֋�*�6�-�"܊o+��8{�]ekC&�N�C1c�¬������S/�r���b8`��(�[Z�A�2���l�ܪj���e'��1����p��@2e��Ss\( #r����i\�,�TR�q��9$�ԑ�.�o->|��u�R���&=P�v�ڤ_>CD�"F���J��/2��ouU
k}j�d_�Ȭ�-��`t�eު���y��#����f�M����Z��-�?PR�ϐ�"�$�~9�B���\V�O��:m�z��|�`��D*��ʍ��ྎv�?T�����4�j�,"��-�${����.�����n�{�7w�:���&> �5� �*�r�j�'�(�m��{��#^bo�TM��!�`�������|�K9���쑶]DW�r//>p{����0.�w������՛�`΁` d��p@��� ���!��ڜx��|�>���m)�)�,GK�_C}}hi,�������D��+6��J�Vp( �?<��N�{ ̲���ģ;���w%C�	���~T�4����>�i��w�J�2r�4���!�����h��D��6�����U5��v��hJ�_u�:�\r�=�\�ܼ��}Ĥ��_�x�Oo8��D���ط��JF��d�̟�	,�� ~�/V�V�K�NF ��nyd�mq�rˮ��T��@������qu��l�O��������!&%�&[ 	��A�EXn��;�Z(��%;�/%yCX`IXfT��H""�|��	����'P���]��ﷴ4���ؽ�OoO��z�0L���9$#� [C�����5���A��W�ڞ;���DH��)��>n�%2�`�ZlY��~e��D���>`0�̨ +Ĉ^{X��� Q��(T�4�κlva����MC�I;կ�~,�lv
��G�j������RlQ��Ϧ>e�.!^�	Pp��{�k~���k�3�.�:SB��!�q��{�+���aJF�5�pw�#+�.6�<8�e��cF&LH��	��[�����`��棊q�Z5���ɤ",S�8q0���e���D8g�8E׍�}*h.
��u����Ȝ���Iq�9
L�өe�us_��I�ʉ�h�+��৙�H�t�����b��M��N
��C7�����s�LЇ%��X�o
�?�s�U�$�-LhX��P$�s��ak�E���#Q�����n�E���O+B���J�vQ;���%\Y�[�Xa!��H�C]޲���{.�x���J\q��i�[�*B�ç�l�]�P�EM�,Ҧ	���J��	G��=)((� Y=G�m�_�F�:g\T��~*<������6e��-���f@�Pv�,g=���	���R�e�CS+�ed5�hH��\�a�]!��`g�vp�,/>�@���T80pzz���%�� ��~�֍��{�����<��@�C��1�FWj�Ă��#.��Au4�9�v{0����[-���BC�H�s+�����M33^e`�m(#����:��D0�Bn1؝���l����T"2b��ݽ�����5��������r�xF����)�{��c`����R
򒟲g��V+�Є��\� ɂ�+�'��y3���/�J2����m-��lCAz�s99i},�ubΝ�����Ey��:�4L�^k�Gd�x�@�A����qf�7�KV����sZ���,4�q���lf����h(V��L�K<�P��؄��ܟ�α;�'V+���ѢE.hFQ8r���g ���S%�;����y���v�]����9�/��kf��I6��=�驇!�n��"������w���>E"��[��������O,��j_��|�H/QU�8}^h�ؗ��[����%/�J5X���Z�ްO�숕���'�����
e��������8�ʨ�4�:�a��\��8<�)����wAI�z7_�n��\W�����2(�����3I+�dcy�$6�*����������`Y�q����9��f:HV��9��I\�ԗ*CƎ�fs!�t�v�0�eR�p����&s�,[��� /�Jd����*"�E7P�T�N����dq&��@�{���7�!˶Ѫ��6�A`��r>c�"��*<�p�������p|�9��!6(��p�[�đf�uJ��3�wO������H��?�l�$�)���xT�.�=PZc�\���Mi�E���3�}F����7���~L,ʮ���^�H�Xʕ��d�/��L;dÏƽJL�>\G{� � ����)��G{��?	7����M�w ��^���D�M^g�[.|��wu����3�!3�)�M��f��˨�e�@��������b��2��b�&�2Uvh�۷�i�>X����(�7M={;�{�W
0ef�CZ�1��o�)�9��M�K�9`�b�]=�5Ǜ���T�,�"��������q�Ѓ��9e`9����.�JD�=S�B�/I�,(���_�y)��[�A2-���4C{7=��RD� s!Z.�ȣԈ �<�Ξ���<�'����,(b���4�DmE��KY��O�&��������Q�t}����CQ{{������L��d���{T5U��S�.L���?�r$;D�~�������q����N|�b�l���v�y|�|�f�煴f�����e�`��}��rw]21x����x;ؿDU���R���q?���|�{;`.l����k�HTG*�q��Y$�gkd��q|�����ヾ؜�hD�zY�n4$\�������b~x���h?�>�d�"E��,�L�D�M �zq��a�'�O\,��������?]�b��1s�(��3ϰ�X�.�g��D,>_(���{|KV�YTƘ�Qiu�����ń�~�r�-���<��oy�HU;L~כ��>�f�V'�mc�`�;�7����B����տ��!l�X3
�V]�ap��W� �v�B��Ts����l�7�����uOPO� �d�����	��A<����a�$��D�<������y��؈aa;>�� -I:m���w�v�]�]gQ� ^&ͻ�l=�,L���PJ,<��K���~x�)�!�����&��u��26DUpe�ExO�ˡ
I�ʚ�G��k��q| 4��y�����ٽ��-b����"����bE�E���J�{�0�\{k�d����H�Os����3� 5�a���q�;L��~8p}�6�0�?:�v2Z��%W�n�u�LF�;�<�m��tr��m:���Ę �L��Vȧ��J?�������\�{9O�{�J�5ˏh�T�u0��B `�Pk��M:�N����(�J���_f�q��觌�.���η�.T�W��oq�N�8�6�,}�B�����Y���j�b�XĦҺ����?!k�JO�c�b��w�<�P�*\҈�D�P�wG�z��Z#�dC��A���Q+;���筳��;��T��y|��� Iۡ"�"CE��j3!P�f�7.����z"��x�dQ�7s��n��~�=�g����u����{�<����gFf�B)�~!~����㾽��[/P�)*��~�Dq	��a�� >���W
[-��T��u.�����~W��-���8�+x?g��%5�����wtt0���]k���>�+�����:�|S��^��L�j�`�L�{%�ҥ����tl�V�۶m۶m;�ضٱm���̜����B]u�u�z����%�Ҫ��Q�����Јa�:�o9͢���M�+Hk�χS�ou�A���P�������J�k������y�M�u��#;�Ǆ��L��1q�t
����Q���+��6T ��:J��3u�>`��yTx��Y�l{"J��A��-q��B���N"{w�!��l6���ixI@o2Ʉ�.�➤�:~����G��ѺueA�(c>I���L�dBOHu�҈'�ŬOeP�l�Od@h4RAP��.�T�R�@�M:�{xF�U���pY$��忴iXw~�U��<��������i�=��[�]je�4�I�D��+�Z��u#����Tsd\�yج}����ڄ7�v�:�T+Q��d݁�T�Y�o�-�!ѽm$ȡ8|�EQ�EIJbc �N�>�I�p!�P	��ǜ��L�Ω~�����4�hx]�tf��#�)�g�p��}uj� M��R�79�Թ�O��&Jb�M�7��I��:�5~�⍶�m�QbP������PaN��].�-c���y�L O����*-��(6..j~YE U�.ߙv;��7���.j��i��3Q�e�����9Y�j%�+0����Դ���������<'��J�5�d�N�K�g(=w�s_ʢ.{f��#{wn�3]{���g6b��?Q����~qFz>��K�+�48���iq���me�}D�KR�k�ЦFj�!����oT3�>�*׆�.0?�_�UA���Z��0b�\/�UVRw�3�8�g0�U�5�7� ��\���������S��"�P;$�	S3iǈ��V�o�X��K�'9�3��0U��rBk���z�q�<�0�)�<e�0mU�i\�3�͒:목�^�9������`Y���'katGx�8x^�N���h,!e�+���r����R�*�����iց���z�J(E�YY�O@1�%+���d�5������=)�I�XzT6ȔN�?Vj�N�W�
^��[s[�l���J��aw����X�Q9���g��7�a�<q�&̬����[�8�]�R�AeP��|ggW���HTƒ'S)�@X�B�?Ψ���Z-��;HŒ�ӠT%�\"(�ω#�d��.oL���Mz���xmm\֥׵���l����N�˖3"$"aRA��_��m�$�6��>
��9Q���K 3D���v�W���.���-���pp(��k[��� s]�My���˺����S&��CkK�D�?�~�"덦� /H���(��X?D0��^��4~��]��em��XHο#Ty��	h��,�r���˿��z��p���L^�y�t�
�z'�GWtD����3q��Ř8��G�mB�H��~�`�b�M��זq�T�D͘P}N�o<Ύ{n�����(?�0N���T���K0�!{z�Z�;����w��@�,�#b:ti	����M���,�U�NVÞeU�
�/�Ï6���kXČr�,p3�aKp���|k�+ވmB~�7; Q+U�P+P�Ձ"3m����@"�R���M�����I�[$�j����<T�ui��r���J�W��Z89=�᝼[���l� e��}G,�?��Wr�3���b�?ߩ��-��KzzP�xuZ���L|~���� L��g�~b�Օ��>\5��~�H��;�d��M�PP���k� sr�����R��N���t���y}VMI�WZH����3_�� \�>??9��~_����H��k����4�Y����g���{إ¡F,�m���ǓKo+~�����#��tBݛ�\#��~��;9���A� ��4�*�y��������_��5˅^��z��	R�\P6�o]Uk�Gt��Ő�2���kwV�b{�A8	��-��f���*Պ�1d2N�8���[����I:zԆI`��m��z�D8�#�Ӆ�
֞`"�P�d9Ԇw3���m��;153rq�Czao�Si��9�vhDlM�d�X�ߧ9�#�K�-��<-����H�[[���󤻛h�wr\E��Op���Ɇ����}�P��P����;�1g1"��` Շ�����m;��WFnZ��8F��8��4|���|WW&��ʲA)E���,B�����Jz"����ڰ���e�<@�C	��
�yhM���}��Ѥ,���.���&b-�h�c�0Ϋ�ɬܜ����GK�?�<��.�p�U[d�Cק�*z�l爠�dko_��B� ���4d�O]7} L�%@E`��'R8߹9�4�l^�);�Ԃ�Z*��.�F ?)@�+��`�ѯx��񱻴b�
��a��1����]9����}_�����}[re������{���	�6þ��v��:3����q�����q�{�svq�d���}��{��YVoR�����?нJ��m�����k���9����=��t�����'4Ҝ�OoݶRx�x�l�>ܷF
��O�Xg1�̽hH�3(�`�x�i�����a�+��a�F��&rR�:�2�i�
H���!Wx9ל�N}߻�(7]��,'w/��tcd;TБ�_��r�33Ɇ�s%L��N�jvo]���HoV�ގ[8?���gf2Vy��5�
9������km���՛�c�F^�*��:� �*!! (��	�w#O���R/-^ըX��A��Y��w�#s1B^�$���[ǌ�~s��q�-� ��@�~E\L��w
��Þ�g�JU�Zwܟ�O-��6)j������ �r@�� �ց��� :J��T5)��,���&{<�>猘O����J�YB]^�SY��\ol߈X����.-�8���~�������h��,,��^��A�r�<e�" ��$���R���^+1.0N��g�X�l!|A<6��Wتiz"!�61�B�`LG��v��=�8)��A�	[>V�굃�x�هF�4�!د�P���X�u6�ܕ��#E�Ŧ�<��߉ZXp�i�����^;��w���� =�����x�Q.e������JJ�l���ǙL�0ɽ�g�1��n�B��j	;2�^�[&�bX�;@a�n>Oq���z#z�g��gR�g!^s/KȂ�'|mQ��^F����������OZ��k�-:�"�m
4E��Q6*D۫�H��&�mi�[��˽l�X\�B��g��+m����:��?��o�Ob��D*�|*���za�?�~XX����{����9�X\z������Pʋδ�=-s#�^� Lm�O���U�n��'��a�*r���#��S�w�`N,��w�Q�ŘSظPg�@kVyϕ��GV�T�����hhdC���e��_ H��ALAQ�SG�&�I���]$(>�k�Ռ��YMhx�j�Sv�t?��i��2��Zjry;��<�-	���_'֩K���~.��ΰh�����Z� -��
�@�]dr8�efN�l��W��B�9����L��:��#ϋ"ʽMW�V� Z�x�v�*BdJ�1�ϫ��N���.]f������*g�����Ms:�Fxҩ8�w~Ru��P��U���_~=�hii��s���x^�)b��Q���T-<���|m����@�;yY*�<C��0wGgkX��.ݝ	�oY�})�b���4��)��a�}�?r��&s����Y�Y9|�m�J�/���Rc%<\l�.zj���GJ�����)�M�°������ƧPf�����H�����0>K�$�d��Qkfof��f~7��� }g��8�˜�����-H��lW����m���rJ��T�r����98TD��m�x!˝]t-����e-Y_��gF�H�Q�X�VM8��5]���i�2�oяʤ|T�G��-z�(�%�bY��=���1/c��R�9c[�G9���p1F�	(H�˰�]<�X;���8_���=O
��c�"�	N��Q=�&0��Q�@(Z����)20D�H�r�^
���Ւ��٭���<�w�
㦖˶���H�X��*)��BƆs4 ��[R|�+�Jj��]ʭrSp�a�4��w�캒sM��4X��I�?xҮ׹�=�N��jX������p���#%���b��8����N�����@Ӿ�BܹC?T���� <G��NiX�MB0�V��qӮ�u)�>Q�c`�=�2�د��Qy-A�&�RB�}�Xl��g�?.�[ˉ�dh���	Q:^�-��k�O���f���N/ls�1"�(��>��}�}��F3��}�\\|�'���B��\��Zm�{��`5]��
D��2j��`�Þ������@��g�?~�cQW�fg಼ ���@��ńT扒��^�%ؚ�gJ��Ն8��fv!��/�l�����8��}��F�϶�g�dG����1�NԔ>��#���P����jrɜ!���#��������T""t$��`���8~q��Ȁ 
�D�����AI�6��ڕ��l��4��G��ڑ0u�*z6ZP�"3@-��!X�~�p�#K�����U#8Ir�&e���M��z�+G�s���B'Nrt�a���i��U�����f�<��2j]��S���HVpb-l(���_$�Y���r29)�ae2@T�o;(�&����Te���h�=h	Zz(6~?Yi�����;1
��y#F-8J:� ��Y˫�q���N $�5߶��(�EJF$�$D&���N%�i���zI�ލ����*�XP`6X���ʻ '=����z笌����PF�����A�V����pQ�T��J�獸�F�q�*�6w�	GAQ���N���~(s���6v���"�Z����np"�7�4��#������l��93�K]D�#�����Q�Ԓ�P�<2V��}�d,�gd)��R_�i�Qw#�w�Q�?��y\b0\Tt+���Ca6̨�%k��x��V[����i�<�����Ʉ͙�6��b�����A������t��p(ռỳz����Az�7���1�F`�?�?EL�k��c�i�`�s�Y`c��)�L��D�I��vw.�7Ũ[�7�:\����A*���Ť��\�v������+�;b�m��&DCF�5t�hY �)��by����ЯQ[ITʅ�yh�-�0��WsQx�#CY���r|��-�=Y��k��G07T
{� ��q_ܯ[z����~2�4��T ��B��B; �QR��00��P���!C���jB���[XP���BBj����n8�hnq[��΍��v����� ��ʬX��c���G�%\�UE|�9�T�q��1��2��ο�oz��yh�ڃ,4O��=������#L;Ɩ�'l1?������ρ�����<M�o��4pᐕDTJŬ���E���e��X2�����������d�y�80�3q$������$%^��yup�ϭ���c�l,3h�B�Ԅ����GN�߳C�)w��q��5l'�<�:A!dH,���\�m���7��s~ G���W'� wv���P�:����HuB���H�+�B���i:�/����O6=*k��G3D�Z�ޤ�<}V�q�|Yn9�65GH��~��}vb��42���W��ܠ	�0��<,�n������G�DH�fFx�@���S����;d���]��F��m׎��yS�E�#T��*�
03�t����b?G0�EE���@i7U��B�P��4_��d�U�Y�䈯8�7:WP�wu��_��s,ƀ&s;¢�ŃTd<�)����H��7������p^��4��������l�5��P�K�M���'�+��@dmC"�o������VK�5]���X=%귦��A�?Gv���+c�����1�&�]�<|�j�T�·�F�d�dbK�g��Ra����E�5aT&�T.&�r�` �(|���-�\	�H���v���Z�"�<G��{�����%�p�7���=
�A���l��;�ص穄:�j.�ku�i:�����`�k�e�t'���$���nb��h�W�ث���e&bx͂E�"�]��q���cg����{H��n		�̉���m�Rb�� o���҆��ɦ�7(((�G�ؓq�d�;я���<#��]萳̅��RJ�_�W{#H��#F�����U�1�a���R���;�Mx���5��Hf~���:k50�r�W�X>��X~��a"Ecq��ɏ���=	�O>�����'3���ބ�3�O�/�ؓt,�'6�_GT�W4���{m���Y8���{f ��d���y���Dv_/�9R�YsV�jx �3ݩyEW�@ ��'�JLo���5T���T/����9�8���g�^��-���3Y ���:�p���j�d0MTwR�������0Y��C�Ia��s������D�o�s����N��`����/���ƣ�����Ȟ�ǉJN?[f#�&���x��3YX~��	����9wdW��MU7��v�0���O����I�ή�HE�%�5T#}�ѵ�|ώ�=�A�Qy���y��d��(���݁��h��W�B���8<����s��й��S�Ӣ�Z�Uu�׹9����l �v���o���@:�,���]r@�����c�ڞ��6}X�}YD����}/��V=X0�Ÿ�9��R�mZ>���}v��@����u�so�}"���,�7���n�#)���K��	�I��VRE3?R�{d�_������I�y�Z�����)�O����������T�� k��I(��5�e�D��h�5d��EK��⏚�Kk[AW1L2���Uc�� �h�i�x���9u����#�:��)���BQ���qlD9�D=S4� ���f���:�KK��x�v4�����O�۾}|PFS���%�9s�׬ږ�a)R�;!�y�T��[K��	[�M*a�U�f��*tư5,���8�'j;���t��ɱ���:HcR�r,����-��2!ᝏ�>�CcV��޾�4�	E9����^���1XL��J",�.rO��x�q�M? �O��|�\B+��P�M:6�%�bЃ�TT�c�eM��܋tP1F�ߣA7=� M`a
 B#
|Eϑ*����a35��)���[��ڔ�K�[�E��7B$G�rE0F����=�\��nL���)L��kK��%�Y;�~��esbFVWV��n�aI�4�v'����e�1'��Fa�Ho�ޭ�*%I���{��dbc	��q�֗A8omm�����G��9ǡ�'pם^�k����1@T�XI�L]�Tb����������9��3D�ӳ��ܶ9��Q>H~��y���
0�%�<�d�2.7���9���V�lam9�7ȩ�IDz�!	��w:�,��#F�#op��Z�%~�%�/OeKp.�<#6Q�����}��ik+��E�K��B�2n,
����\�J������b��VB�����ͮ�޼��A
0$�l|ʃ{k�Gլ�J3` ��*՟�&ks���`d����ٗLn�:.�c�apPD�p���z�4�p�,�5�©�l}5��v��hB ���"phd�HJT��~\�n�T$��_�2f��ZN�3��p��8�i�����~���(�oT(e�$+Xf�s����X1�laW�A�JY�8����pW�&]�������0��I�?�KtD+�OBEm�cVB��ǙQ=�[%>�oA���X$�6�����Ǹ���>���E�ťZ-�JC�',u%��q��N�J�u(�*�A���M��^�zᩑp\l�5ɋ:v���Z;������������X��@8b�8�L.�ڈ�`�1sb*�c�1��>8���p���%������Ǜ�M܏�����K�"$���s�Sm�]pe{�aa-~}ZV?x\Ջ���;x�������F@D�/˶Ĵ��ܾD"��?;J2m���;���W0���m����n��</Amp���� ��j1܌�h%��3�iEA��G&36L�9Tq��
/���}� ��E�ퟁеvMQk4��-����%�ax"F����ҳ;w�]^W$�0��9Q�ACTx;∟Y�f��J*�� ?)����\��_�8�ф��c��R`E"�c%"�Z�!g:�Ad�
��Σ�*N=5����~��o���ic��SR+�ST���� 4&�>����ـ�_hh��k�Og�u_������Y)%�i�6�"0����@���Y���a�$.T�!q��H�#P� @���h�%�	�g�S�!�� ��C��d�0�.���
��Р+��e��C#E��'�J)��`#])�Ja�>���}P�Ȃ*\�˻����\���N+=���:�䉪{���8�,��=��_ �F������m?����m�)�h�.��[U<>�\$�[�U��JHsO���~�L��gœ�&/)i�#�k��G�=#�>�ly�$����y�H��gp�)?ٗ?q\���*��T��e��[`��C<ܾ�
c��'��0��s��/��11�������;��B�%����{3�vwq��c~�Hس�+�t[v˾��[��=��<�J���M&��[�?>n�`�@���r��0灮$��nܡ����͌,��&�̄�e��
-C�S��L�L+}�fdq��+?��+Z����J���l��C�|�F�b����s�,'�{)�_���m�t��将-��HNT��9�7"Zݍ��
{^S�x?Ӵ�%��	ZZ��d�|��&!���uհܐ��ֹ߻��>�-.�~d�KA� EQg4���V�)�%�Wf�q���ݖ��f;n��F����JX"��+���.���&G�����a��=��E)47�Dĝ�r,���M��)��U`L:pti�"4D�$$tYU?�|{)������� �<ڹ�iB�L%�R����JD��\�s�8�-�6heqĺ��_����3¯���������3.���\�RJD���A\�xT��������c��.|�[Y��X��:��)�Q#��I�(�+Gw0����k��p��<���0�rsΦ,'�D}w����g��Z�Rx�p��|ĝt$)�'�Ӊ��4�7��
m��f	�|�[(i��S� �%[[H�vok����kw7|�?����_��X���X�5���o��M���:>�#�ǌv�Ր,G<��3R���f
4�̿���{��� �D?�3��	�.O����oMx�7Z��j?���a�r=�1u{�+�����~�湭B�Y(�tܦ�`B��[�0 �K��7�V��@gJ�+���M�������8�v�Z����լ+����:R c� Z��#��/s�t ,��Y�� �����`@�ي�L��IW��|1	�X�✞@�<�p��h�hin$q~mԣ;���ގm��C��:Ԏt@�@�yDg-2���޼�����p3�4���h�f�[Q����h7Ҋ�TU�F�|�2Zf+:D��TD�gr��]J:�M�����j��W��,>�䮮6�]������gҧ�vRjB�/���|����x�c�׍;1�on���E�����38%l�Ylff՛�M.���?k�Ǩ�r�о�h����R���ʺ򃚎��Y���%(�*�LI�A�<#�w$�XQ{���6�ڳf�﹤؂�K�:-)�c{
�|�b�`MS�.�&�8�������������������{�/ub��#���#q�-�X��!��p��tɳ����z���O���c?�_��&=y_��Afe$��Y6�	�!�,@����%6�<�(7Pw��y���W��9h3�w����[�Hw�w2��.��{Ô�~������^���Q��Ur�is|��T�J0E)�"O�j�GÊМͺ>Eh?*r�~S��9Z@�$�hp⍥����ӝY����*ƀO�1�v	����ڡTz�����[�qi���,$���w?�M���$ڱ�1�#)2k�LgVFq��R3���@
����`�S�z��#���F����߯����6F	���:$�7�����N�(��GFcC�v*_�I�N��K@�?��?�Q�6�n��?�N
<���lJ�\���91��%��d㩅�G9P3ˏ��)<���y(�$�~CASI7xk$_�t E�ҭ2��UJ�; ���C@�TЬ���U������@�Y�c�o�y�*�n��/K�E�f�m�c+G�FU�]X�74��/�:}r�vW��AOn|�i�߇R��z��s��7hs�;\��u|ٵU�*���YʏgZ�"��%��v-��T{�f~ЊBcm~߻��Σ3du�;�+#��_��5��G_�b�o��#�����v5%��<�Y[��i7`��B�ðB�dp�����+��.���:ʈժ���fM�X ���^��oG�{o`E�j=�����)���J�~�>OR-�DN�/�o��JP�g�.\fY������Ʈ�)�g�fjf#Y�_��>ma����&�Km?�}P�mc�3�W��9��J�u5�S-�9��T�fkQ���j}A(IT���5�AڊG�J�'.x��ގ����u\�A�r-|( dm-��~�z�������{����M3�)0Ӫ�do:�9sb~ZZ���>�h��L�0�4)K��gj~�����<����U{�HI��Z���fы��������m�>��u}'��R�dDʦs�`Q�G�}Grk�����#$J�Tu�-�]�_uw��Ғ�oN��nn�?��.`>���e���"8���rF�_�=�n�+��pe��5�[}��L���{C��d��$���(,��"J9������ު�f#�3#��^i�Vw��ěp(19�����K0*����$�'!�F5�t�+����c�q7��~�O{������y�#�����w2FLq�w��	��I��!;�����9�]o�pqm&J�؛�}�;r^�?kB��WO9�àםi��[^�w��<�MDQs�$�\��1��;Xs��[f��iV�'ۀ��_�{C�y��0F ���OYH� �Ga�;���U{��ݶ�����5�?Ȩ��l�4��s��={�6)$$�wvѮ���M�Q�>:?���v3p�Y��}�Y���#9H%��eY�D��=^#����uѤ����T�uD^l�����Wr��T�"�x�y-��'���*�"zR�Y�Q���qP�zW�m_z�GR �N4,�$�s�ʱ�>&`_�+��<Z����8?�VK�,8Ip���΅�J��WS��c��a�����H$Cs?�u��	��0MsE�B����*(w��*ǃO���7#��.E�Y�E�v�_b=t:v1�e��p�C���-�>���,���[<��X�|�"��r�&����8J��@`8j�_~x�^��ר+� /▗�[R���Š+�QK@�_Z՝?#KS
�ygy׳�m'RnqV�@'>�v���т�@|��	~�����J�����p9�
��I>���Mp�a�:^07��v6�������P7�0۲p�}��g,%ف��;��iХIMv��~/�|�*�FY�pxl�'�X~p�i�sC�sv������d��M`Ō��,�W���d�F-b���eL�:-VЯCB�bY�����wc/�嬡�S�E]]0[���x��q��
u���@�@p�Z,�Ɗ���&��?�����x/N;v����JȆs��b�m���të���X��7��E;o�[+�V�eP*d���V{�Tg��G�k�,�8�<E��'.@����LL󑄟��T��?e)�b �"Eؿ��s_�?�J��o��+���6J]6�EE8��.t��2��DT��zNs�ȩ�c��fK��nZa�΂zoa�j�%N�BlA�<%�AnN�S	������<v�0Ӻa������p�x �hȈ�!%1��Ǣ��� E����ȍ������	�(V��<X;/S��� �x1F���-�8�Ji�w�Y.X�-��}�/4�O��[;X���x�E�C��M�xEJ��~�a
��9����l�J<���>!즃��������:6�>lLMj�0��"��_��0:�,�}��)v7~��>݁���[H��������H~�v`���7D;,/c��n������ d�M�8�!�y��I_�GN1��dyqʽ��bm���}�1ۿ��XUUB�K.�7�z�+P9Č����5��7[y� '��وq��/B��Nf��i�U&C#k� �a���.X�Y�[��"ı��W��8�3�'�?�*%_P~�Tu��c�
L�+�U����	D�q�3Q�����ʤU�yT-UY�̢|��㟫���K]�>����Ͷ����Tq;A���������y��p���ى91�}|��_�+����s&|�J��C�Ч�NVN���GB�O4G�m�յ�x��T���t��t@O�ֻO5��g>��\nVv����, s{�M����E&���y��ϥ ����#��g�]�v15*���l3a���e�:��v�t�ze1{�h��<��'B�6��I�1��[0���r���O��"�i��_��DO��\q�!R�L����(���̈́�TG�M����x�7�銆Xȝ���򆳨�b�}�Y�`v���r!Q���Qf3�5D�!�*e�,����yUy;X�������c�-�|>� ��[tWB�ā�z~�����!�Ʀ���
����������p8Z��C,:y�D(�o�C�nx�v��A�����[�tL��p1���ى�
E��E�B�H2rH�1j�p����jA9�"���WD��¬,B�$ʴHR{��{�
)�u*�K�4�R%D�t��&�,�GB20R�ߛ�;sX���^z�07�{�O	��� �˻8Z-�C���k�-G�q�Jw0I���[�[FM�{�z�t/|B��6���֊�&�U7��{����T�>�^ؕ$\Luڴ��{'��q��?E<���ɧ�u��l�|[1O]�/Λo���J׹�A}������VG�W���_6��,������k�2j5B�aΈ��Q$@�;W��ڜ�H"�������l��5Ϥ���p�׌	O�/CA�=�J�J8�d=��yE�"A�F>SNeq��+Јv�s�ܑ��뤪0�'˂�53�xsdA����i	`F�R^��j�Y��ʋ6�h���;#pԑ�pG���	��/8@�z£j��C�WSyQ��!��L:�G�esj�1��~������̀EZ�6%ZëzUg�s�mL[WR/�C��RC�����~��~P�qXD�����~k
��|D���$$�� �k�
�{�u,M�#D ]i����lRuI�Dy��ڷF��	 w�HabDB�tX��3ҡ~_��u����%_$XQ�iK?H�@,S;y3�f���2�P2?��A�������k� s���5�� 5t�e.�0�{Z�㳚_U�j��i\x�al��89�5��qA5˃���+*0�H~��d�iY�-N�ј�����pJg����=���z|��htR�$�������K���e���oo��f*����ClE�MN$E�sR�~�i��hBt����B�����!�̫w��d�����)-�[����+����%�H1�Ms�(�]1�J��!+�������i��,آ����3�7�����g�P�� `��|AX��f"	q�2!��QmaZ���!�S�"Y��6+u��q �4�+�����q�@4-�9Y�"�h���ӱ�rȸ"�U�z�sU64�B�:����s9�,�����+h㲝�	xP���-�鰃��q4�4�({�+�t;�V�Yc���N@!.�)3��^4�D�<fŭG#��1�nz��4��Gҽ��bx
lt��YX]��*O����V;��Ng(Xa�2v���3�}�� ��^9NB�#�To�U�5zG�����ws�&@�S�6����7�j>s��pl�򦑭\������[B�����w<��	H�.Z뀅)�t���R�Y�	@��IZg鐽5}*���n��K��﷼Y�/��^��kH��Q�<��ϲ �o ����Up��њ���
U���Ð�A&5V���)�&O���$���݁��E&�����hni���h˚f��l���X%�=���I��HK�N̿�(�:2����'7�tP�7Ds���#[��z5����E��q!�i��6E$b����JF� ��\�8�C�t�HK��U3R�`�� ������@8��	�x=SU��:�;Ì*؞5n!�ddN�>�B�'��n��\�Mګ\d�J��-2 ��[���� E�Ys��®j|�N�	x8�Ā끡���ŠR�t��9������~IZ���q*|n�͛�ߜ�|���UhL`,��r?3:��@�gɨ��I'���'鋔��XH#F0���\�(FvK.uT�HH|Z�D%+9�O��}���NH����3L����xq��e�dX����p�2�2T��� 8�iŘqV�t6�0 :��m��2(����d&�l�^~_E���0g��\ɰ��,]��,�-�'��F���M��&�����9����&A]qe��K�:�����+�kiF��覆W�Y�faj��ջV�OaF$��'���B��5�l��]��W����)�[�>�X�����k7��Q���=�<�u��� �ɴ��H��k�r�e�P
QVg���D��gXzNBc��3�~�ך�ն7'�}c�O �a��"��Im0������_��+`���l����7�5�CKJq��m�z��ZA���[X�~�����4&�b���l�X���^�K���>BJ��k��ul�q?�����e�Łaۭ�/� b�����	�.�o@b��RSw�	�,�!��5�K��dP�A4g�,dP�A�v�Ȟ���e-�]4�A�6����,9�a{�i�u8/č)%à8��/�:�M��_&�6�B�v�'3�/�L���z���}�?xM��&i�[�V0��l���H �)���27�����	9�;~��n��K�A��}^22jR%5�F:+""$s�(�	0!!;:r�[�����t�6�Y6���ƿ���b��D��u8	v��*��Da��a�?�'�B8�bu�c����Z���yn?� #�gg��B�Dz�2��x@m�����{����U�H��>��2c>̄\G���j��4W��!��Ȱ��=�j}���&���l����9�F��,J4�B�Rr2%�L�Ux��|rE�u���$�l����ݓ��Z��[@|��eg����:�7���G���J�7��%PL��^3�8�q���e���n!�Ⱥ�a��OyV�L�rω�q"}*8�c����m���1Q�`c,�O�N���D6�<_C1q��J�9�.�Κ�кT.���6�i�T�V'a!��G�ݗͦg�V�n^(���D@&Ym6ӕ���ۭhq?�ݲó[kurx �ܒ��I �)�;�e�{R ���Z���h��3d�䬂��u=���9$�t��$6�8�
Ez��Gtwf�TslV�R 
!z�đ{6F��,����0���6��n4��yQ���ㅿىJ�Ϊ�v;��q{���w{��R|���S�\ɘy�4��It>.�d�u4J��(����U#$t@�򺫑����ù�{ʼ��R'D�BNXteA���yt�v��|0z������Y�):͵�e󼨯9�9g�%`>2�>���C�dЏ	w�p���.n�tHdZrH��O^0ɓ�%�Z�Wb��|"���C}��B���j
� �J�'��3��L#QФVKB 3oh�g�"1&/�%����fvt"��<eڶ��M����#VB]3���g֐�,c�g�+�����9�Yi+u�� ]���(K�cVg9��J��yDd�ũ*�/�����&]H�E�i�N��=4 �:�XQ�*Ͻy�HJlg���)�ԀEp�N+���DƮK�l������Ǚ��מ<�4=�TɮEv�'3����h���:��~��}S~d��㴝���h�\����/�;la�,�u�psu�d��5��xaZG��V���s�PM���1��6��qp=Ŋ\܀.U^#N����_�dO�=9�{��kF�U~~�����]��t��o��~�ʊiN�j \y�F�
��K�gw����b��+��%�sb�vǶ�tl�c۶m�fǶmwlk�;�>3�?��jջjo�.Ȝ;��ڃ�$C�3fH��~���hs��M&3�=����J�GF?����:a���-����p9b�o��<Ҩ^-�UK���eFj���M�Q��l9����������Ӕ�a�٨2ސq�;`�(��T���"" ���'�����s��mDx��#Y/$EA�Wi��!7�O��	Ф�'�!3�
5����֥�]�LEҡ� J�£�BY����q�V:�l%�Q��׌��W��27�������O1�Ǣ�LUu��=:�]'s�PE߯��F��=/���ʭ'6R� `�,*�3��\�c�; Y��:�1��'���Pc枤��E&V��B+ʪ��8~�����/p����|>�E�p��b-�B��������8�ȷ/���酠�p*8ЇCΟ�޾��(;ߗ2w��fW���B� e�j��o͝������"?���^bd؎�R�'��j�A��l�-��GSJ��^���x�*RTYH�45���pa�8���^
C��Iz�LaE�]w7��k�]Q�S�+؆��d���l,�$,	��j�<f�5�u�����7-���r,#`��Tf��!ڀ,Z��_���鵁\,�9P�"-6T$���#�$_�[��N�R�O{2E,3�R/�=}����-'MtS{ш��45D�8v�-�9�h@hi�u��`��z&I���!B�Z5v��h�A��B]k8���.�S��%O�A�+p$AUD��IZ��x���������sw�'�%�,V�<�	�Vu���k0Wig�rA�'
������f�����y�3�f�2�<�@�z��%��!5��1o�r	�L��]�f�{���5�X(����@�(��&�F��'f��ȥ$�ڣ��1f��?�b���d�~�/⠦�w��q�Y�$Co��ܨЃ5��U�E]7޺5B�7�n�0�N���o^(���d��8ń3�)��i������ap��i�z�)�t�ol������,3�+r69,������Q��U����:�UEPH��+��Q2d�1�\�j,��ae���`��G���.�u\�{�_V���g���wJ���( Mb�����h�*ճ��9��^���!�gH���d��V����:4+�vx	�^�%�L?��ӄ�ϊ�*�GE�!���Y[
D�i�����Y~�"����>��}
)t(C��Y����O0 $�"�!D�eYSB��y0G�� �[��ucS+��L�=��ō�2�w�l������d����]uR
�zi�y��g:�:t���w��x�7�;L_5�͇3u,`���4�4��&H��p*�!�j�E�H�P�$��0HÐY*�}����w9pZہ��}T2v���NJy�4%^3u�\����դ��Y�T��;1�{�V�
�`hd���J���d�ܹv���Wv�	��E w^s�~[Jo"{�q��a��e����H�aX��q<M��*q�DG4\ywpk�W�s	��r"3��Y'ކ�(34 �2;��h-v����^Hu,��v��o�;1����p��^	�k+1����
�t�_j=����I/�υ�/KLSR<����p�HQJ�$�,;�1N��.�:�=�H#wP�s/��|�n�]O,��3��[��rv4�'����0��c�j���5���F!I���}�-�h.]�<�����:|�[��*����uϢL"���p*��П0Ȉ9���������`g�������������{�V��{~�v�٠�]��6�G�-�"�����V��M�Rwb�����<^��8��/ߧ�����6��x��K��@�ǡ��*Gx��]�:>���İ���_����j�Z��s���F�0�^�����������r[y��8~*+���}�,,L $�A���_3��Y�ԏ^l!ĥ�N����"����@��LZ��p����}ް�Ϳ�}q;����-r:ɾ��S]ջٱ�cDE�_�wD����j0��6�z�Z*�'c*Xq����l�}�f����`bLO0�g3ɅJ�NO�XG��=��9�A�ԓ������6�]̤�ڌ��Ͼq��U�����i6�±�t��k5z�<c.�z�P�`C�k��	᛽�0���ji�5^A��S*�L�=�m����b��Bt�l��@QRo��!��I���S�D��g𧫽�y��n0��܀�f13�jZ�=��q=��{��`Ӊ�e&���5wy�!ٓ�`��m' �4�5p�:��>&u՛>@d�'ra* +`%�0�N�	���<N+hVI��[/�>M�����:���������r�3�@����y���!0�9LC�������v�Ҿ_�����Џ�wy�P�?[��h���z�����}��s�	���I�MQ�u	���|�r[��6�K�*7����o �B�$�i�նՎ��f���w���+Μ��E6�� ��5Ox�����N�o�3�l�)����{�ǢStÈ���#;�}�D�O�'re�t��a���ğ<���N�}P��O�ف��.�x^�͙{�ՠ�^W�׺��)ۛ>��.���7\C�����ϪKN�B傌��������r�H�7�*�Q�_�V?
�ݤN^(NH��pա���8,�����%I6��P���o͟ ��m!���|� }Oߢm�f(r��i��B0X�Su��we�6G04?]�0I�jl�"t*8����4�'V��z�h��/U�4����vqnV�_�PKf�i�֬CR�\>�J��7�6A!��$�J�܂�CLl@�����D�Ȩ������C��3��w�uk,�j��]�W5�Z�2y���{Q���hc���\�{3]�7'�b�y
������iO�����J�Ϯ���emxO�*��#h�(�Mr�30�x3�I0r�	�\B�A�<���WGđ;�hc�{ܢ�Wk`n�ımz��O��@"������c�D�~б��a��
�[1�	���Q�.;�`h�Mh���j������G7q:tԉ5����BW��{�Rբ� ӕt��zW1��R�3^|W�~�QcQ��%��2�NL�<�:�i)�nV)�iBCu���5:t��ggm��w;��J����G�P��ߡ
�S�1�g��F�Ǡ��gBo��3wG?W��	�a��ʵ��~٣�_��h��^��C}8w��s���+����n:���x�*j��:_V-M��#�,�����|>ly��qH��KJ��s%��tԺ��dk���*�Ѓ�u�(�<�9WזD�UL��1x5��q0��Y���Q��-7P��ob��(���ꕒe��O�z��Kh���.����ʂ�n|��(N;����B�<0v?�ېS���r14�1�ۏ�]�
	�+�M���Y�w'�
��[�(�un_�e��:����(�Xd>Q;����K�t����A�U�>>v���w�k�\����V��=�ә$��pq��cch�<+U��_�>%��:h�`a�d$�M���~��D;�Ba���/�6��8�OީND������ؼY��d�ZZ4d���$I�5�
NK�!qBh ��q�0�E&�xxg���т�_�O���w@S�@Q	e����CW�v�Xʥ�����da�`��d�a��aB���0��Y��O����Y�	k`�R]��IX�ڸI��~eB�(��k���
x)oϥ{����F���Y��l�x�W���Z���N2	v<B(�j�rN�0����.r!M`-<�����᭺����|�O���j,���h��Ե��p�\D!`�w>o�b�>���͜a��q��w�i�#?���tV�ѫ4)o�E3��@3�9)��!|k1$�M5_�4�ێ�pl�k�ɠ����mX���B�c��pD+6���X�0SA6�4A�'C�����:��!UE��˒��U�6�q[�<e7wu/D��;vȖ�w��u�oD�2W�SD�wZ5-/ل�#�P�3���'gs�h��Ft��t�&5������"ɉŏ!Vt\��)y�U�'��L�h.ש3�s} 7��k����&k�v��![|��w[`SJ��M �*UيP��kWw�s��%~N��c�QqQ�`����7lzL���*"�L���X-�s��F��GlV� �YFE�GR���雜�*4��y8캽�Q�P+���31ԗ(�J6�$Nk�-@���ύ	����T�?�>�P=3Dj|�R�0D����m�e�����(;��j�[DY˲ņ��`r����w3�[��n�Q�d9�-v��d�}�����Z�{ke�-���t�����QQ�8��/�*���ٻ��#/&�{�n�ن��R�]��L	���݆n}��%X�@���j6o�q�;���,��%|P��X �U+�E�>��Hu>v�'��S�h�M�Τ����ߨ��2TUqs�m{���%q:�r.�Ý�I��A��FO���U(����]����kN6D@N~� ����8T|��׾��?��']M�ùQ��F"��k��ڰ�L����7�
}�{Y5\�,�V�>{}}��d��~���BI�X~4<������\ɚ�]ʟ��[3E_f�Z���NM�kZ:=�9�*k��t�ܡ�C�Ʉ��:Z`&3�aO雱�ǭ[g&�����=��b�^Ȳ�~%��o�E~F6t�?�s�62��M?X��v�iv,�a��!��o�w�,�빧�С�ߟ�� ���m�u�fjtQPC��e��ʈM�G�C7r�b��>#f��3#���`k	E]��ó8�Z0�T?�8�8���ұ���N�/�I����'%�gj
�r����R)G3���h�^�C�, n>c8�/�����䯣)N"9���Jzck
B�*�3\OJ���������.����0��uN2��Q&Z�����=��4m�lG��c'F�1-�|c-z#w�؏�Ve���Ƈ�7))�CJ��OYw�I��X��W*
��w��za9���� �Q8�=���|�*��s���i�,������u&w�BdD����&K�.(EFN�~�������;��r�e�'SǄ�A2���-2n'.Ǯ�H�C2���e˳؃h���fߔy�Ƙ[2E��L��\1�V�ɒ4=����'m���
.:b��z�=�Z�5Ҹ9q���7<�E�S�x�~翤��yۂ��r��1�ڥT�۵_�CK�4�v���$�ռ���9s�jr�eg�Gδ�b���P����,;��׫�ѥQ�]���<���k�_&[A^~��\h��}d	}�^/����d��-2�H�t}/�BiUƑ#_��/������cf���~,��?�!J�g*:�.
<��03c�(�it��Ֆ�Q�^�j�r�܂,#`( Vr��u�$������z�;���O̎W��,�}��L�<x�M=������.���w�VtE���Cf��z�u�"i�qw��L k�܌2������oG��;��L~t����|�l�!�n�~&.��j��G9HG��Wk�S��|�K���3�u�!��v�͜�~v�k�rc1�&��#L�ﴕ�p���զ�n7ba��t�ּ!*cCsc��0�J��W�㮎��Z���3Xz��T���7Q�Q���BUsLv���CJ%�3�V��p T�z��2���܉�g6X�UgѨ��l3���Y�q��N��uFY{�Gg������7�?@�G�FI#}f�&�6M߳���K^��.�E�UnV�*�J�=�#����Ӭ��{�e�1��)Z�x��������e���Yچ���Yg��@
�q�Ab�I�oa�.<-�=�����M����"�/�s����0��BN�
z(�p�!,v����n��Ր�V���$�"'W���������Z��a�#h4yu���(�l>�V�����'�4�OV�YA���R�BR�6�b��>$�Q�M�w�N�(s��4�o�'4ێ3i����h���z|�#nFR�&��t�h�����m�4;��ͻ��	,����
�7�HS FMi����f\�<擧���=,�jJF��=��m�Y,z�._h�?�c��e�Y�a���[�����Q��/͗�V�o�X	�p�8W]�[���ߊ��Bm��Z���{U*�{����x�E͛j�D<���?�`�o^x� VT��}���,|r oe�D��ȩ����%��s$�V΁ە��K5KW%��⫒����5�-,��ŵ9?#T��ju5_E�HF�-�k��ơl�I��1t�ll"R��d��`>â_��.�i�����CK��#����u��n�ږ�]�YF(���RU�Ώ=$E�;�k�WU9ټA"����)4�W?%��'��7��S�8af�cdh���|as`OC���HH;������~�ˁ?��{2�%q���b�5lZ�4�h�ŧ���y�6��	���� �A(=J?5+u8_Kn���� �������#�b���V߮"��a�O�G��C<�M��+N8�8ʅ���CwU�"I���m�V�e}G�\�TD��L]�Q��^�9%�h �p�� %����� AŮ)���^W�J

F���?��u/[�Sw�a�ݝj�r������ 2:Ӓ��o�
4���.��$�A�Q��]���VR�
Ѩm׍^��x/��2i�e�5ʳ��Oq�L�]�,Q����Z�y��OY�I�vb��QK���&��`�hs����$ͧ�P�ń �|F��$�ႁ8�A(<ã��v�ߡ4I��2$͓��lu��l0)�J%�;,^��J���u�KE�M<U�D��P�Ɋ_ѳ۬�ҝ�2y���j�h��W{>��!W�B� yĭ�m8�7W��f֗��X2�}{{Pϼ�h|��Qu�oQ��B�Zi���w&�z><�P5��l�M$�bG�''_CCLrE<��ױq�S��*�O�H�Ѭ9ԓ�P���M��+U��������odbS���%ɠ0��a5�����r�����V�[��B�*
�e�O���D뒲2��*Y^�W�?X2�� ۍ4��A �Zt�G�v�ɉ�1V��i�qȹ�����1\�\\?�o���Gsžr�Б$�[S�*8��d͙�/w"A!sՑ���o�h������Yf�o2,-囂�������Kf���Y��=J"T�?r��ka����GT�x%(Ԥ򫌤Ԇ�9l�/�?��ד���F�z�u=�ś��ȊM�:�a��ǂ:��F���t`&)��5̥�_eh<����'%۝�������UV&�O������C<;��o/�=��{�C ��;漦p�A��D�]m~��"<:�r��d�'��V�$�*5hͶ�����/�EwʉIOe� !ʽ�J#�R<t��嫵9b;�NUw�-\|��\
W�:��?�ϒ�t	�n|>^�����]��S�*ń��Cm�-tG�����!�b��:ԫψ_����A@�%<��!�J��/^X�ɧ�)���w�������e�[Ƅ2U�Kӝ#�u�5$`�>����"q��2�����C��Ι��� �eS��I6 �5~�W �tg̀�Գ}=lt�㥞�j� 5A�;��y�s�@�5�,�sw�O��p(���'�Ɏ���|)����H�@�*>ޕVctg�L�߸Q��5�l.?�C�h��kF�#a�5��s*W��5�]zI)H�㶄Ŀ>�Y��ȫ��Î�B�M��`���Ш�\�I�3 Cj��?ƿ���(ݧ��SV�ނ>�|����hj��<+u�K�3�|��2�������cI���E�����:�g�����ߣ]Gc����jy_��v��γ�
�7�R���4E2��hT���������1~^��d^�:�6RB����I]u� �yeK5z4��eٙ�C#ư(6&��(�����%�9ǦF���uY���?-X&�Gw���G�z�9�2���A���8�J�H�Y`<�ܼ�$k�yr�ل�P0���,-�̯2���T��·���L��v%�z��� !aq������̓�؟o�ˇ6����T�ëo��3�<R�K@�Џ�EQ��ssF�?⌌C�\DC��!�,G���'���NNN��ď��y�<���R��}^�Zw��|��^/���4�@F�8Iv�im(� �/ۦ&Ģ��?�q���j�B��뜄^�܉�m���7�ϐŠF;h�����u�73���q�QC���sq 8Ȝ!�~�V�����}��W�Ek&�/GT�܈-��mԛ%�\�v�9��KS�*�M�#�󓏢+K�O�q��T���'	V��+ֹl��T��c��T�����w��1�(i
��_Qۅb��)M�0�#�J��_O���mX,��?dM?����,�<j{uDd����UAnr�������$� x��g����9�5��Ԩ�M9�ib_�ӥy T9kv�������i,]*��+�dv�Z�j�:�d���-��������[��}b0m�??8���ۍ^���3Ep��Ɠ����@���S���+1�=!�R}�	g2sӅgSE͍��z/t{#s0���z�8��~>=���)���~����h����N������i�B�N�Ch��nny�m�A�W��5���7-Λ��Bv�
�'o�L#�v�߶lC�Z;��
]��z�Ol�O�@^���caŉ�y�K�T��#���m�������Գ����!;d7�Ba�6�����i���<��-?mԡ"������H_�?�ڶ��M� �tb��?C՟4u�0��P�f?���`�Nnܨ$@e ���P��԰�:�Ȭd���J�[D��L���?,?�7��)����������I�����;=8��7���P+��E5�Zi�z�=z2�x�x����U�&��A#���`)ܴ�r u���T=M��g #��M[�%���&q6/[�[Ɉ�n�� *��е}�UR�¢SA{�x���㒪.�س*�.��1�m�P�i�j����I�§ߙ���Bq#��� ��
�\1��;�FJ��V?�ѤU����T��7K08�F����L4�Te#9�ꐪ.l�Y����Ԗ7��h�P�����$r����W���k���=�#pg��)4�D*m��EO*9]8.��O���� �vV}��ߚ��O���v9胈��_�R&$?�tv��a�	U�K�5l4/4!�8[���ª6���k���|�q����š4��~���0�� /�U�c ]�H�!+���l� }8i]�M��Yo�	�z*_�a�vLM8� ���"�$���g�Q����J_��aeQ�K�7����6��]�5�Zf��-�(���Ҹߔ��SFII�v�T�>���/�ۄ&DF�|"��l���#{��@�GW8&J���Z.n��xJ��lL,2��ƞY�T��_?N;���j7x��x�`�m�4⼂8`r�#�
C����q�ݮ�������+�B�~�g+�>�ףĸ^����[c�XWO��*��(����mU	ٮgw�;Y�f�k8�b��'ۡ�q�KPY߄�`I3�j%��U��X����\J�l	[U��6�e>��%������I��b�9P^�J�5�����	O��*�K��Fn}K�A�G����o��&�3�R�B��K@"����"��l�񯛅'4՛� �j�Y�e�ϡŪI��H��(?�o�g�i��.)�5�3u.��r����7��	���QEj�����E�3��X�*F^4�]Ѫ����<�7�σ�?�n�>��?0������kB��������\Z��Y)h�ɧ^�ߺ1� '���������U(�E�F�x���fBN3iNV��9ު���f��z(K���\�D䋨�d724DfQ��`IɅIф�U9� 	��v�)��v�FE}�{�"�w��iT������x������N�c�2�}$k�j����/�1Q�]ӏR��yM3�5�A�e��T������iNM�dݿ�F�0�`vKӶ�CO�o/�"B�k��*�'h&�gކ�\��6x�%6X)��HO{/���坏/If]՝b�p��"&A���~1��B�5a��Rc�|��IGp����!�f��$SZi\�J���e*�
t�ZpօioiP�ç�_�ÀZ�e�A}�G�YOA�6��ܨ�����\2:{�G�zXLj ���#���`<�Ȋ�3�EF�`�4?���LI�D�D�j���8����ծ�e�0<ab��y'����CK���dt��yŒ-��pZ2��u�N��$y������C���|κ!��h�4��-;�ԭ����ҕVQ@��BD����U��w���$/K7q����%�Pmb!���V4�%���ۀ��"���f�{%�ĝ�p�6Ǽ3 ,b��?�ܡ�&�\�M�q�W� ����}��\~	�����h��/�G}`�K�ש�C'!lM�k�"�ި��+��()�ͬ�?��DCI*�o[T��lUV�㗖s�"����&���	(E3ƽ�[Q����(J�0S��/7��n�_H���+ϡ�.w�� �|�'_'V{cաۉҊٜ�eԭj8�j����?]�}�'E�5����]u�g�ԑ�ҋr�q����Պf�=�ig��Dծ��94縒e���M�(ol�GQ�SV3��h;x���p�i
O4��/�"t���y1G�P�hN�:���1'�(�}L�A�&�&�C6H�+�ʇ���U~o�:��e�[�&F�6�M��hj�v'�3Y�_K���&�/u�Zc������B��rU�Gk�M8�b�-����z~�О�+	6&�J�	YF�+���a.�d��>��Y��n�~��u���~#P}�@�ܨ�kNu�M�?r�
�1$���j��2��8�����ķ�ʄ6E�h}z9�J�>n�Z?d���+;=��_�!�D�~(���_*��{�ة=�>]�J���x���sH��u�ׯ9��g��)��a��4<}q7�'ǜ;�x �� E��#��Y>~0��3�Pt�� .�Y8+b�KwD�O�rY����:��@|��9�I�7#�9� i%���ɗ*��+��vgMK��8mť�Cf����ZO�p���SF�O�"�%2!�E��-��$-ab\-G�o#��%��R�������|+i�*m�kZ<\S������/��x�y���g�F��Y���-Sӓ�[tFL��:P�;�=���P�l�$CO��Q�}���p�īN�]�y��$f�4զhJ*+�-ɫus$�s��I��i�91"�I��߰Dm`�H{�t�yޣYư3�q�t�d��d��!�[�L��}���}2��gD�&�M���X++��Y�92���
?d�ENR���h�*^�󢪼:a�:y*	J�<�b0�Cm�Yo5�DP�s
Q2y��o&���%�����UU��83Fr��)�|��t�A@�%�"�KLu&�G�����%4VR��7#~1���^3�F�MV�"��{*���Dm��s�9	���B�U�G���8..�î����T\p��VA�O���<�t=Gk��$��c��g;)�oS!�""!�]��|2�pxI?��7��a'?@�� o���[�BM�J}(�����g؋��E=�7]�WjU<�&W$]\	b �&�+H�/:I��R������L�il>�V�5�>��s���$Y��ȡ,QVb�׻�p����?L}2M���\"�4�+t��^(�`iN�kQ)VZI�Y63J�1FZ5H�:K��$�_P���.���r�#�E~�L�V�V�?=�!�R|(�3
���u
�J�>��q���K��׍�uZ~Eȯr:n;�>���1B?�8<Ohi {e��%3�z�xN�\G�gS���ʑ�̦+ix��@c���`��p���ͮ����=&D�����4xBvI&5Y�8��}���o���Y�i�h��?�m�\��V0Rn�M�b�#S+��ڷes:dhj(CLY�f=|����|�I�{� ��W81~�a1 !ʚFe ��R�?ʈ�o�o��N�MW����c�t��`5��bp%��[��nw�ya�7�z�*�lTW��)�#W�;|�Qz�\�:F(G��X�B��ڳyE%�u�(!3�JM��r�xAO&�����#�$>8��s�}0QҬ�oB=��qa17b*G��+�����tpѰ!��W0���,d�i'��pUdNЋ�[D�VE�{,����h���ۯ�|+��I\��"��"b�?���\�&�Nle}���v��R��w(ɠ1�:�Q�Զʲ��t��&�]ݲ�r������������5���O��7��I��Io*�,�����'�v�;��)���]ZN��}�6|Af�����;Jn��
�%�5��L�"V��H��p�
�lΥU�"5 u���caKbF��{�C��m�5��}�u��kfZ��J1�_����Ks�3��pGf���8��2��T�	}gwǂ�q[���6be�9�W���F��j���Y�FQT@+�
��l�ӏ�ɒ��Oت��""������F̳לٵs����S�5jK��9��R��~�Q�P���;��x/��!EI�Ȉ�C7��Ɏ8 �yS����qE�Po(�#��$O��|�J]��ƥ�.�®�X��&pWk���x<�JY&_�����4,D�,�n߾ i��]]�/�n��GF|�]�R���&p���]5�ޭ6���cn�[��t|��I���7Q�&�eG�qHD�4/�����8�-5:�����u�-��y�IsD&q]!�t��~��:z�2��v{�7E@Sswh�ʨrjy'p�*|���,Fl�H����荒�h)l����sv�U�Lmsq���I���x��������
��l(̸Jf\��YV��9��D ��2�I��}b�ȍm���Z�p�&�y��"HTu����b?4^Me*�úJA�Š)�6%o����	�-Y��� �W\���в��6LAN��i=�Oq�Y_N��Q_;�H�OX�@'�|�ث�sǞXnĈ�Uʛ*r|&��z8���~��a4�`C7��!�;��D�{�r-خ|�ji���BNv;���;�z��%����������O0f����,�h��w��)w�m�n �J�E���bs�7�?|LK�i�Y=�B�Z�tvD��=+8^t
��e�谦�b�zST���L���6�R2Ƞ%��&`���Ɠ���d������ꪮEQ�h̩��yˀ)-� �B =tV�1��<�V�-8jg.� ���2��X�ԁ}��[[���v\��I��t*!����d|̽qfX-"L�$QK��4G�!�Y{Ξlw���̍��	D�'�)YA�Oè?&N�ɏJ�7ݑ3_'r6
� �48w��͋ړ�������:�;to)7��1׬�4�|�W�~��"���G�<p�!ͩ�[���;���H^F~�$����n��l�E�gj�w�G#G��я�{_�W ��u�;���7u
S쁁�x�K���[�)���1�/*H�a%��;?�3s�p۴�^|/����-e�ϋ�M�ɉ}����������0����[���W��2���D�"�>����}����cbDU�r�Bd��Ј��-�y��Z��Z��a����[��9�Z9�Ҭ�W��s��㼸l�����O.���������y�'0��,V�h���Α�*���f륏T���;Azw�A� o��VF�#=u���BH+#f���~�����V�M�J�����S��4��}�m��x��z�]<�o�"�}Bny>�+Z�Y~j>IY��s���/u�EB�&�V`�mܟ�"��J�`�h'�\6�3��g�j�W�)߿K���}E��ނ��F����ey�u�SX�<��� 1��dNz�̆]+��g������'��9|I`��ţ)��VK�*��xQ�]ܪ�9�^+L9F�GG�`���ת��<�R��R�۱�:@\>v���%YV6+B�P�kS��qJ2��F�>I���鼋�S),�yGXO(i����5;�q�i�̔�`A<>�,I��Qf�Y����ekNeA�87SZ��:���R�l��eȪ? ��r�;\�N,e蛴�����.�(��CD�I)�?����XE��J�ZvP��ƴ(u�Z������t���58�C]��3ʬ"{��,��A�����i���!"ZZsu?���T�Bf�(���U�'����Fv�2׋�j ��H =�[����~:�O�o���d���ؑ�/XN���C�c;ܞ`WF�Տ
�e�ܼ�5�ei�	^��^�@L�V]_= �q�Q*	��o�7�{&h �f"�4�����	I#�"�-i�xv���u�ʺ�@��Л.�@���E�泗�(@��ro�l�(�� S7"o��J,C��-�"J�;t`d%q0�Ȅ�{D$R� ^K/l
�E,��L�������W3��T
�3|�5��sdj���e�4�+*�������z�c=Č�}��Yf�1//)J���a1���gŲq���uM~+�D������6H�H2�A���R��j���B��7�5i��� 1h<�R%m�F}�x���f��죧��O��k�r��7����ND繳tPn��_w���7�˽w�ٯ6�EƇ���#ɚW�����(X���!HA�:��5�6���h�|�c����\W� �h�x|?�k�{)u-_���ϼM=2ü)�0��$V����}�"���s�=g�G$R��2M3$փz�ie�	ÐrG�(Iq<G��F��u��v�i�����! R?3��Ě�E4A6�zo�<f}(��L�Җd䔙Sǽ].{Ҕ��w���ΝQUZ�
��N����z�������X5�B����7�ZKmj���˃3o@۶p&�A�=��?�&n�lH��v����bn�N��)禚F�g�{��H�}m����Z�f ��+��d��{wI�yH�O�5%M4#�G�j�]�腚��	2o݉�
������0���D_���m~�Ѻ���4�6(�1��\�m���Z��fQ<!_%a�K�_����Ǜ����jT¤�>7�$����tK>����-��v��L~L�tI����cz��8�%ӆ��H�((#-������VAF�XY�ǃ'-�:�����C�r�D�8-8�6�C��q����sFw��A&<QêE+����B}���<Bm����m
��Bx���"�x-M�ec��5�|w���;��8St݆�/����K��,߬Ug�9��k��d�����oZ�I�,��`.Δ��k��r�c*�6с~t���O��v<I�(�4'���U��������L̅�tA8� :����N]|!��O�V��i�3&��07q��k8�0��z��7�+r�l�99��b�G���譻xF�$O�c�rlF)~>}�Y��F���B�Qy�~���IN�*�`$i�bLG�a�0�1[�IWB��e�{�g����@u~O�	I���oϑs�?�?����*��&�<T�h�^���O��S�X3����;2<��yx����c�C�l��*���1g/���zލlY
6Z$��G�r؁�qf8}��n�D��&Y����w= [��Fg~�n���ؑ�~��{�8�
�r�S��U+B�Bxu�R�d��Ce���B�kն�G��3N��&����^�#?�`�.@�M�Wr���@v�������\��Jz)U��H����$*�bIA�.��4"���of`y,�S{Z�)-3��9k<�z�J}�3��u�ZY����E��֎cC���/'l�8n���ѥ��`�gji)4�U%6O��/����=ܑ��}����%j|�0�N6�0���mEߋ���U�-�L4�Q5[�stq򱅕���i�؁���7b�UXu�:�#���1õD�Nⱄ͓����Ȉ���Wq�%iS=�Ԗ�#VL���LkU�$xyڂ5ۢ��l��hW7�ܞ�:]5�N�c[t�����J�ǳ]�'�\&�4�y��lǿ�U�m�����M�˛�qRk}Si�ZF�_I��h��[��L�cL�2(BɁ���q#�][H�[Q�ۻ�������L��-,��Z�~�20y{tj���}�Vl���狎,Ђ A�l�N�GR������݁-��ޮ'۶m�v�\'۶m�u�m۶urO<��߼3��;���{��P;�)�>f�L��#�dmO�wi􌲈�i]� ���04D�����'���F`6H�����p��5
��NM�O�P8�"qkW �E\�D4��~� �ɧŧ�宰ݤ�]��I��:�����-m�>1�-��=�F��$�?�,�8��oH��s�O U�Y��b^��|00#Ҿ�$�BO�"�:H�����y�X?��������\�F��PvU�=�W�b�;KŧL���Y�����J�
�|s"Ӱ�`��B��F�� r���N��Hܥ��Ho��h�wCJbh��
�n�"x�ժ/�D6X�S��>��>2�جU�!�R��t!�y�_�m��N�ێ�M���Y��VIN0R�K��=9�O*I��� ��Gm��tK�������v ��	V��Z�ᣑ�cI��Hy��<s�2mǎ0%������Q|�����0�D�Pf`K���e�Vڱ%��v�	���)���	���ҙ3{���Cx��<6���"-�j�b�F��7�ˤU���26�d]�Z���e�t�<}{�r�������،�W�k�|4�3%z��G>��̴�+��	�v�/rg����og�D�,A�!��aY6_�����GQY'[�=,y�?���~�+g)%��5�����v�Ew�xf�{�pN�u�Os6l��P�D��+�+�̚pd���0%�kk��� ,G<���J�!Tc�f�n�MK�6K�����ab#���Pؤ+I��	O]�����d���ķ��}~5 `55
NȘ����J�o2����ˋ�|x_EM<��3&��]O�B�
o����.#14}~����2M)ML���Oڣz*�$���o�rk&+W/�vB�4�������Xu�!�Am�!:0�껙��Gf虓gV&}��H�׫WZ��2'}�"5��!����B�����)�i�����LF�Ĝ��S�C`E���WO���'[��m�<��%-"[#�UR�W�nEh�B���"-��᩵��*�rGX�#HW`��{�{��w�����d�y�q���/	o��B=p����_L�l�*�m�l-{gm�Q+�Sb/�X�7۪#x5�{�.���Z����l밥*�'˙/�Xnr�����'�ԛ��oy���+�~+0z%�yC�:���O�g=��J-���=W?�n�A+	� ߋk̲o��AGǅ��E�fk�����hF��4��ԛ��m��!�^�,�%a򗬛~��M����:�`�ᩯO/�O�����U&_"�泾ܲ�9��r�W,�/�J�_�"J��5y��4�o�9�N8N����8H�6�o�}��|�Ă-�ON�"Jb�5c��?ٌ�����\Qy�'���F�nѨ�P���\��꙰����E���˝�ku�1b�����r����l�t�uu�j�����wk�=���8.���Bt�#׭��婳���WҾ��C_�f�t��.�ťҬ����,Cc���
��ŋ�ɴǽ�yh-������E�K�_m	j!e��W����jC6���l�'�=�n\F�Ag�5Lt����������y�kU��|�|�j���jY���by�GS@h�3���ԊJ��jC:d�8ם@w�F�b)�8�=u�l�T�����&���m�d�t(���t�@�SD����'�f�$�O`�Hqn�c)Я!�{/�fתFm!PHF�θo1��(�e�X7ș����+33��mq'C�e�e:NR!]ۏ'Ŕ�R�M#�\η?�nCm��H�E�_:�q���~uAdH$(J��H��ge278��m.;��h��j\�3���{$��Gvx���v��ݐ[L�6����o��!�shP_�;�*�Nߜ?�޸+�t��ikfV���o%��؛ב����%�A�*�9�7�:w�ɇ��XXB7߬�����L�3��i��mJ���6�������$��f�UY�/�=ڼD���'y��1�ˁ�!����:�~uwc��	=��F�<��MMD�F�y�� ��V��p�Uf`��y�6�B�ZI��� �߉���s,r%���Wi��0yH����}���$U[�N�$s:s�PM�
YX��%��D-�P�E�FҪU�r(pU�����R\��Pk$��)��	Y�P;�D���*��+��n�=��ԅ-�uc'�ϴt�Yg��T`���c����n릀h}��m�qi���Ŝ�I�@���{\n.w`�F�-c�LJ�1��C�^9��渞h�:�:�Y}��	�}��2z��;̋E����b��w��k��	%$�20��mz�v�>��.rӯ�J����?�㎗��Z�ֿ~�9e�r>�n1t�q��#Bw�hҎ-����J�˩�ƔaTK÷�V!�WM��i'�Gx�CXr��w˒Ev��Zu *�u���1ba;t�L�!jt�����l�)�/�DC���n�5g	&�������	(�����L�Q0LI�cm��a�]uǊ�J�ׁ��f\9 ےO�>�iRj��y�[&nM�7�2����\F\_��z:��e���%�?��&��HrDh�U�p_�-i+�T �qQ��)��3o*���g���(��].��E ��� ?X؈<DY9�w��w�|u���;�6�ɦ���uq�����
l�,S�%&�������ﲲ+Ŏ�eD1�����4���p��0��������JO�@	�<���d]D������>��_Z��D ��$����U�����Q��U�s�CQ�BXte��s�TRW��.EG�ϭ�[b;pp��Gi�z.%�ma��1���N3Ln����V�)H�u�F�~
�D�:�w��&'�����7�~���%n�z|ˣ�+w�������7�m�$�ˠ��[Ma�:A��,���|�{}S:��"�"�! %?S��wDޕ�m���'ߜD�:���F����}�q���4^��׈F�B����w����)���:���ج�CX����,6�Bˈ�hL��\ǜ���Q�ls�#���B��n�r�3�v4ㆣ�m���lC�
��
�
H-fy��/x��<ƳhG��C?���Q��%��B��j�9���5K�)�lΓܻME����8�^��;}�v�V��d����̙� �HUWƴ��wU,i��D.�F����D�E Z�DA�泤Z�kɲdogp�@��IK������zlG`�8y�&mXc����~��|>V��~ ������Mz�a���*;��&8������+�l(���l49!�xG�M[��A<��N���%��'(��u���w�CFDD��aw&��q��:t�l���Q�V!��ƥ�jň��f���D�IB̐��+�U�%g�@�z�Zp�[�r\�����`�UN��_Ƈ��3��˱��(![^T�3`��� -�F�cX��[��}f\��W*��O*j}�F�U/T=��}�cC%R~�ٲ3�(( T������i��-:��T2Q�6o�7u������gc�����ĕ8k�R��O{�㻟��D��t��s;��/�{vl��w	<���8�̫]����"��G�C�7�*�S����#������u���C;��g�/UVE�^��5mP�@nXq�޼HW�����r�GFehӥ��.�z:$�~��;?�N3p�����x����;�hkH�ƹ7��+�Ju"P�p�|�����E��G�����8Z΃X@����~�Əaآ�oksK1�b���f�_^n��,L�}5����F�N<�2웂� ��.�m�S�I��1��_T�%�P�۷���������"=������s�Yx�8��))���t
����#�Y�\Y����,�����k�/x�12%��<�+���?�s3(2?sǀ���~w�G؇����0��~_���?`��4 ��������E;[j�EQ�hQ3���w���TM�A�9��>A �7Q���A�(	<�<�cb��㓧�ʰZS�d@����d���A"͟*ѻ� ��D�B���m�ZG�"������r�b�&��E���7��, ?;X��Fa�]�Vxc���P��X�+I|a�	��\t����w5yg<��Y��93b��#�{!���/�)�a#L0��W�������;t�Z�6�Bu@�5�!wH?��`?�z�N���9�K��<U�S[��� C�<�IV�pZu��S��D��q'p���̴�y�0Ί4����Ra�Ñ#E�q7����z9�́8P!2�VT��3y̞��8҉�%?v�f��e�O��GW������ݶ�c\�	Jp�b����.F�LVH�/�L���h��R��ܢ^��+�jf>__�ŕ5~h���E^�ыFV2�Ŕ.���n3Ù��mj>�V$�-xU�kےv ��1عGkv�S��9��Z~��.e.ܘ��`�8����L3P n�\:)e����<.���f��^j�r���y�D�t~>}�m�P�?���p�F��Q���q-bzB���Ck����t�9u� S���_uܟ��ic�W��&��C+��>V4��<v��4����p��:F��|�2�S��dȊ�~�?0��*غLH'���1[�3���yPn���p)jr�I��c�P�|�o[������6��BF�_I������lk0����G�Eı�9�7o�pd�mʪ)�p0�UѐG�;�e��kt��y_�b��q9l�+΋��!cFPu�4��dK�2�$`L6�uy���5��(�����e��+I#0�LF%Z�����\$;����{�R�bc@�
'�+�T��G�Y�SBVn̸��CIF�ֿ�U��ZE|�����.-��H���R5��L��W={�{�!�w����j��Cӡd��c4,0>HX*�u��h!]����u}�3��#,���4��g��ē�$�'�Od���9���Ci�Zo1Fp1��tT;�٘F�Ax���H�26�̎��ڢ?���z|y��\ac&����O��̗XN��G�8֗Aa�5�̌ ��I6��	����M��{Y��n�"%ؒ�����.��6^������R3I�g��S��>����s�����,�(;�7����!��s���Z��=J��+�7r�.	���c�-����c���p~�A�d��&Z�����˱��CQT���	r��<�(���k�H��+���A�?����by�|F�������$0�V0��J�k��V���IZ b%�ջ#s�u�4y��)!�`�V��=^�ݲ��z�0����<)y�
�c�*� 9݈���0y�"���P�v���9Ė���A��w�
���7��K��T����/kB�P�7Ht�Xb+.L���ay�����K�n�CU�Կ0�����A�����-y&�	�em�˳��y�������̣���}�[���(���u�U��͸Z����?�""�ôaF��c�%�L��&���	�ӽEW/q��B!�=�������+�Ivc�b���܃2�ttt�2�r�]@BC�4������zKf����d��7ۍ���8��p	�7	�Z��E��(k�>]d��l��Ģb������pZc+I;X�ya8O+9�<}�/\Ր�`��\��s�h�q�� J�r�*"�8��y��g)Y-3)W��K?�}l�j�bF��oo�^L��T[i�$&ڙ�EQ�9�@e���y���K.���#i�_N3�k��h�C��2������#�c��	�nd}b㞢��D����גm����B;k��nb?}%I��c>�[l�����z5jISdI�[W^�sA��A���sX+H�@�>Q���� i���$�i��Aee�����l֭���^�zت�vJ�WML�A |�"���U���n���'zd��>2����
�h��(�!���wy"�L$@`Z���0\�j����D�0]f��ZRrB��yA�{�ʰ�V�oAٱ���o�	g�Jˉg5�^X!��g���B2Hs�t��R��h0�)\�t���P�J��"���m��A�'�_D�K\�m
��he�"l��J�׳_}�\PN�N�Uԫh���N-:4)�|Q�{��}T]L�JE#��W�_\bd[>V,�9�t��r'�B\k�������,)<޸W��NS���p���Ԝ6?٩�������M�"���D�A��D0��7�^�W��P3��V��@x}H�>��v�O�*b��l�k)dN�{3r�F��E. W`mm�-���v�]֛�˦)l�*P����wC�_�;~e��nő�K,r"5W�;�������6��Q"��QD%�^�B�}���~��_�l֣�
�67����M���3X���W}��0bU'�=$��"�a�����޽Q��%��n�F�d��� �R}zF���\�P�l�*_$�(����t�'��ʙ6�X�bj�Ӧ�'9#N�Ga���e+6vM�;��O�j�� }�hlv�}�@OI}�ijW��B�.v/g�Sgp2d=��L�����/�����%�E]
m��z���Q������}��b��P��,�:;F�T�,�CP�)���.}�w�l5FUzcn�����B���0t؅�.�<�˕L˶]·���n��	�_/��-�؅��C�%e.�Mi�b�Ұ�]������j�5�Dõ�e�5�I�l�/�
�9i���h	�	9/r���!ٓ��^��s|(r�̉�����d�ė?F@��k�j�{����e���=��t�0F����PDʀd9��dQ9�!T�(0p�UlyH���F�&�tvZ��ܽ�=���ծ�9y�0��t������O�G^o�G��@�O��yű��oȼ�������$i�)��:�f#��(���pR�t��!�qЎ����Tʛw=�_ Rh�S�8j�tz�G�<�S蓄�f���ƎeMc�W����o^nG�����Ral�������3h_����V�g�P
9�k�df�܆.׳��p����M@,!�;b;�]���ͩ/�����u�K�ED�y%���w#� �g,�u��D��Ͻ���u�=N���ا�ediI����*���ؘQ�����<}$30�χ�1W�@��)����7���9�K�ep�������
�ؚ�F�;�4.�$'ƙ�U�U2�N�=�&S�tg0
���PrPr�E��hW�N��'���B�3������fd;��d+�O�#�H�
�=r;�a�sf'L��~�ݶX0_�巧=_m]�+��
t�S[��E#�~56�K�xL`�������q��== � Y˻��m�B��mN�����2�z�Љ�a��:#)Jjk��r�"�(���-�Vx�=��������ڇ<O�)_�9�����~�I�����_��
����q_���f%��߂��O�p�o�*~�ީA_�~�,��v
S�'����3ošk�9qЮh�{�m�FN@T����ǥ`<�7�}d�/�N�#���K}��(In}���Y
 �� ���<p�/��G�=p�������)k�Cr=�#�� g���,n(;e^��#�����[ʦ%�0�3n�$�sf3�[�QMU:�LNo�֚����&̆M�2k����cA��(H�?����"�#Z%> ���O�=�k-�>\w�?�L���h�jbA��J�v����9�1�b��v����š�'ʯ)g�O1��J�̏ĚU�+q�,Yޠ���е�V���=��b{�;�����:JF���j0q������a^��e�\�������*�˫L(w�����x��/ �����t�&�Yf��c��� %^�4uɱV=٪��N�|]\�+ZT+�#��@U�V+�737wD]�_!�1�h��Ŝ�MD h!ԯ�j���Ҫ��b�h'�?W5@�\�d�л=��)��tȂaV���,��DVD���#u�E��8F�&��xN<���c�"�O�hl��0�L�P&�x�}�"$�X`r��
SVVy��rr�Kf���G	�Ia�L�._p��17���]�>_�R����8$�T��(s��XЗoq�2��~��3�B�y�]?tzU��dV�I'Lf����0Җ�MSݡB���Ot����ȑ�"�l*��G�^o)()���9�^p�t�Lb]D�8��+h2� �\j9��&�à�C���A�ǜp��f�L56���:Mu4x|���VӒä{^�[��FRdB/ ��Gu��w	��ZYY�q�[ғ��z"6u���W���I��P�d!!z5h����@�,�\/���1��ӂ��X�K�a���f�3���a�F3�7�^�����u�|!�F�t��-��h�3i������+�5�(}��������mL�8;C Y�OՆr�,l��)пRc�3����r�E+ջ8�:"�m'�eȝ�MS�Ϝ��������p@��ڄ�1��q*�$��_fRyƘ`Ne���v�[�2�m�0p����T�h�q�p-6Sc�ϓ���&0ـ"�Y���8�p���&#^�QXpr�s��C�o{6��:nJ`���%����'p�p|��[+���ܙ��ğ �$�.�~+��5�${�W�]g忩ʆ�j����W�#;#xأ�a2)BM(Ѿ��~^'5�P��8z��G��ΌT�9H��uT�������l���	�W��z��g����=Y�<k�0&R�zk���f�o��,��5{��
LS�������
��nZ�C�6�4[�FO0����[���Հ��ܗ.eW ʄY� ${����ݝ�A�H-�R��Z�t�?!h���۸N2��f�Ů��Xΐ���3b2d�M�}Z��-_�\t�H:��ժ�(�����.?"jԟ&ZǕ^���&6������&&�}�%�:����
)e�F�lw�B���M��O� paXB$aEeX����
'W�z}7�ۘ��^�X��9c(J/��'��������ͿnIQU���b�^�����#<͵F6�5�̣��b ��.շ����͚����.�k½]���H��l*�p��ò�u�j}���� �v��Y6'�0�|�X�ZF���k�@�@S�(�QP
 �������^��DU5�8��g�/=[3�<!j)0�����o��z�<�z�Z4��"#oV���TH��R~'۩Y!R��}7�4����@�k�ͤG���޵�ꍖ�'W쭇v�6�ʂ3'��im��pRGv��xS�1G�{5�c1��v��Q�!.w��KY:�;���S=a�^�g��<}G?~AӋ����涊�t��֠K��!/~��q�z�`��(�\m,}��-tLT��]�S��%�E�4g����r�W��s�"q9��yt�*�v -T5Z���,�-��M�Z���h\�����c�c˔RQ�3ʑ��Ln1ׇ�!�x��*���c��}�|T���My� 6�#��wo�NT*!�D��eX6H�<d1{�����)մ�<��03�蟿l\2�M��	?�Lv�����܍���&���i4�m����Ͻ"΋'AW�&�u�P��^��d�"�{��8�Լz.�B�j����s	b=�;�ɚ���}�gD�p�.��3!+���b_���ǋ@҄�E14���d.� Ή��P�Y�t|,�踟����9s��r����Cs������k�o_�x��@<"(�)�(��:E^��Q0����]\�b�ѥY��L�A��Ca�����N=�>�`k�Ʊ��O�L�|�?���ߥ$@�2��N�*����h�����́��\Q��K�lΆG����ȿ,V�5X0����F_��������ꀹ�IS���L�5W�� �GB�u����(#��{����Z�C�	%1
zSpJu�^�FZ��[�a�I�Q~=������#��`����Pb�[������L"><l�F��e��3b�x��]nl����c�w�%ݍ?(�DZ��V����ʪ�^UI�4�н:�0�#j)4D^L����#���|zO63ck�*��|�94���V�o�{�Q���pRB�����l]�������
�V�A2M��-�j�^	�ɉxw�9��3�#9��v|������9R�A�S��w3���蚿��]���������1/�%���=��>�E���0��]^g��l~��2(@L���8,���n��S�#��^W���7V U��d~���''����i��~�:M�����`����&�ݷ��GM���ci�����ס�����E�7;�ց��]��2���������&�8���������y�W��%x_.8���!�G!mOE���UrE+7|eV�vs����c?�3�N�d<��ȧ�e*�6w�~�_�L�(�g۝H��"�����J"v��ie̓�	g,U�)߹���]���Ǚa1k6z���`�4(&}矑2�T!O\P�J�������i5�u[K��_�iy&���0ZCa�%N�,3�b�3�<:�}������L-�w�$��V��[/����q��1�g.x�2Dx�VF���断�6��|��&����Џm�T�H*��v9S��e�Es	�t������kt<"`�(����A7 Inz�-�NG���=:<8H	�%�k�I*�)�1�8����|��N�(7�Ů������ʘ�-�!X)��{�\�����������W���K?�p�4����r��_��lpi�c����o���Vp#M|ŠO��o�n���q�oL]��#"�w��cpl�,^��(1GU2jW�:�1Qs�����G��,����>д%R��Ԗm�R��Φc�G'��>4uB�u��0�������)�q�g�	˖GL���1�S����p�m�:)�!����|�y	!#�s<�~lmy~(��l��[�܏��e����+�;���������%4t���䪟=T�i��$H�����n�:>�j�Y00��U	s_��a+l�ScVv�l7�zu��}�i�\<����c՚�Q�clVp��W�猲��2r ���/��VI�!c+��`K���`VnT��+ ������/��u����V�iR��;��hF|�'m�y_�zQy�0w��=�I/����j6]�r�`�c��{E�����L��� ��<��r��X�~\Iq��j�!�����,�Y�1�E�^�z����?C1�t�������}�ㆮi$�bL���2��+�����]N��7�!�V�V?��k�T�rT���y�33�QN7��rg#��:t�5�p7_-��7׮^��9�f���+ޠg��hU��9g�xUiq����a,���c;Ϩ!h�����C���'ѧj�e+��t�ܳ��Z���̑n�jWK	�1�~y���G,�Ȳ��O�QW��+ۯI�O����we.���<m\'�;m�Z��4�4�)�e��f#��C�nFU;��o�Ǣ$��j�՛P���0��N��p7��`��<�܀�gV�4�YdI�T�1��}�Ё��]{X�5ʃ�l� ��ɲ��3�Lh� �4H����qk�v$�Db�*��k�u�dٹe͌��mre2��������2.�R���m�r���'d3���fv������Ypc�#�~�s����24��'����rOn�ST̜�YYd��8���^� ���	�ͣ�<�#I���>����F�K��b��ЇD����"�r��3�G�?/��uU#������8ѥ��@��[�M��;��<���l��r��µ������9��Bcɺ�p��Ns��k��4[R�����	|8��<;�j�����	{Ŗ��F�p� L���&3��3�	����U�e���|����s�i���g�8y��҆��5�+nY{��{�a�B��Cy�����?�r�a�[�n�Z���;�	z������!9��u��	�����=+30���:_�w�ϧ�� [͵�m����%[�[鱒�w��p��q�
��vpt�e������'.���:�y�ש�s�x��
p�Ɖ����;��¶�FJ/��wxJ����� !�QDm�ӆ�k#^|ρZ� uӱ�̺�2ֈE�쁬�]g>L��ט��`����r̻J%_��0<'�2�GmbâIf�Trcw��^[���(�����_��pnȋ�{�o=H�j����W�W�x�)ϟq��İi��ju�������2�<h�&H���I��Hu��-�1�g���(g�d������ɑߘb�2�1�~�bæ2T#ĬFP���I�**M���%��;�����VjE�b^�6�#ӖZ��b�>�r��D����	���<����F����=�Ɔ���!���uCE��A)�7㮞	����9�)K�'��Qr]�d���4���1�#,ha{�3��Ͼ/,Y��Lz�~m�v�*�L_�?S�,�é(ZO0ν<����1[h4��������r�@�hQ��Pd���+/h4 ���h�7��B+~�r���U^*����\���� @���Ƭ7!��D�F�|�[f��kţo4���l9��<�+m�>��a�bMT�	��=��;|�_q�J���!4*2�_-$�y����[���i�b��=�������<F!_�l4���}�꺎�Vd�'L�}�(���L��I *��s\�A�D��E��Df �!;6���vԶ�
퉓�0������p�'.����v�� �3?�kYn�m�%i��!�ͣ��k���"��Š���_�Tg0����}+��s�N�Y=�*���a���  �O�Or/|�Ogh��+���u��ʾ#!
 R�W�b�����'^LC?�d4���sT� x��1�-��� ̚�8'���4��p����M�Hԏ��5�p����F���t��f������T_A)�D�*~\Kn}y]�.CNw�T�!��
o�[|1��	~�?��^n���~��^�v/���~�}���qeP4+�W��lq_�s�M ���uH��X	�=N�n�{�b��kN�J~&��}�,�w��a/j��[��Ӧja;ݐ%��'�Z�_���$���dH�}f�@ua�����fl�KT�L4��B}��:0a�FQ����d�D̼��	3������K)D�:1�N�"��[�!��*Af�܄��c��9,����<�����C^g�0,��Rw#A;_9��^a��QR�w�������`����, *)���S�V(0�}�(cr�8�
�'�7@�C(�����:��uS���FaQ�W9\b�p�t?L�C�ǿ�R����iօi���Ż��..�Fd�g�4��f-BM&SX�S?$����Hpu-�(/�D8P�e?�p}G�>%A�6��Uw����`�܉��}�E�L��ſ8�֧K@�s%$�s:n��۸����ח����~�eS�j���F��qt��e�ߑ�ŗ����i�&y��Z�dH&��5;&�2���k�F��°}�I���x���=�q�;\r~ ^?����[�����h�����hb�K	�s�>;j�2U"�I������)���K�+Hl
Q\Uv�'L\�M@�~��J�i1�ֲʏ����bg�]��.�lɝ~<��\�Tb፬o�gb�6�<:�_�ɰuа��(L����J�����2��!�Ey��a��Z	�ẕ�a�T�]�w_I_i�e%����^�C�;B�g�.pI�[���ր�52����K)���-�����)����7vl�|���LC�S�-ӈ���{~>��**ҳ�:4�*�M3!��$�i�*���{uWͯ�6w�{�Ψ"qt�$s��Q��>!@��	��B�&��W���S��/�q
���)ӰK}vV��q~>��~�+�}�38}��R��"O3��~�.of&�4y"�P�_��js6�{�����JJ��#=����h�~��c�FS#�L]�������/(��0�'��Q7P�j�@���EJ���]E�ʎ��O����`Wk
G�??��JB��'QZ�j! ��'�����!Ԧ.�f�Tp�Φ�kQq7�D��'��7R��[TF�cN�gXN��J�q�A�p�܌849��7���)�8�=�u��IVݻ�^{���"R9�W��ױ�ܭ�ގ����!ls[���q����nx��%'Kx�Kcb%����Z��o��G��TN{oڶ%�YQUN�X��T�+�:���ѵz�F�v���?�����#��s�)����Mf�%�!�v��ʜ�b�6؜�*��p:�"H��z���T���|~zX�5 4V{լ�L[1+���G�ԵG�jFY�J�4���/��fh&�|Wr�ziΟ�j�~��S���s��_8n�X}��)>�~�
�e�5���;��=5�)W2���bܙӺ_�!֭����)Νъ�"N���FZ�a8�Cf�	Lf��쐼��8�w�P� ����������o1ځ �'p!(� PG�)e_�ʤ��O�����#������U���Q
WJ��ɧ羁`�1��^�#���У�xa�2����$�i�%���rW���W�m%��@أ��iİ,5-z��4�b�ڌ���`��D�9���<���>��C.)hj�)��q����;����-JG���R��Z� �5�ě����q���G�OL�2E��M����+��Yy���w��{+��+t�嬎����0���E��z�Y&1i$*UZ��S��7�9D���DZ��0/Ц�Y�.���1h�0˯�Q�����@�qg����H�Ko�N�U�@�~�}�Jbù_��#��-l�O)�t"=�fx�="1�-GK�~b�X5'X���柸<.̢75�b!;�l`h��&���>	��Ϭ�͊U�?���.i$�!�i�ci��}&�� 	�"���ț(���X��R�q!8[Mڏ�"��|P����]��!_�BF���O�2Q�F'&��U4��e���ĺ:o���N�k��ɡ�;*g��-��(���G�����e˖F�r�e�]�M�<�g|e,���B*^��ˉDv���B*� �/�-��Dqqg��c�� �hZ8���+� ��U�U�2� ��dAd�U0�^z�����B\����RT���%W���uf�:��;.�=!K�ʍ�� i.�ԃkuj�L;��l����o�ɏ�����|������=_����mp�ƗG�H���o��A�<2�3����-p�+[��y�$��ꮰh��8eC��6��c�~t��+����+����6�������76��t�SH�5D�Λ�R��,E�Y�.L�7�4�^K����?�TԆ���42�bdsn���OZx^���:y�S̊c����%i�������	����oݒ�6a�]��:a���͒1߽�d��}�yٌ�8�p{ĺW����@����J9V.��ѽ�H��V��]cr�����GᎨ���R .)��jWW��V��ޓ4�<H�_E�A���8�6'=C̙z�~ңm[Ղ�6o���{������it���:2���Q
����+�Ɨ(��i�f<�|O�|�n�.P�,�Pk�����%��}#�$~�QZ�B�-p����3��d�S�:ë�݊�KI¸"f��R
wVFh�2��B�n��ݳdD3nd�@��a�e�-��O����B����Br��ӯ�)���2� ���8)r[���+a�ڪ��Д�Z
2y��m�S�B���.�����F��aJGf�%�H�!T-6�����˲@��CFڣ0��M��i���Q��Yq�w.���me]jt��u����;���F�l�b�.�FO�g�4tC7 )�^5~F�M��L$���j�C�I�<������<���4��{��GRk8T�1X0���Lэ�m,�p��h�L�~�]()��n�3T2Q
0����H�}���D�����J���O���$N�cJ�k�ֱ��)ՊyvP�W혍��jΒ���~n$�o����I�Z�$���i�H���}��a�qZ�!?H��%Nnvέ4h��[�4t=u�U��K�7���Kf��i^�xE���Zr8�ļ��,mt9ffM�B�?&ށ�h��MVŶm۶m۶m۶���تض+��}�>��z��}�1zFl�>R�e� P_�0YY]'�R�B�.�!/}��U�iue�$�e���=8����} ��H�	�F`1l�$oM���=/������z�I~�p��'(T���Z�Dۚd8~{*����,U���9�'�p�q?<Pw=�h�>	u��eD�6*'�U���DF<��Yy^�?�YP �yNG��QЙ�{�M�C^4N��d;]���?+���4C|�8�#�v;t�r�`�P���*N;⋿�<%J0�����?�^nk� {�?&��R'9y4�d�)�떋<,4����O�&��U ��G�֡�����d$4�
�V�)�R6	�ք%Ӏ�h��(Z-�ȅr�~ ��4�#4��_N�]o)FlDd~����`��h�Ŕ�Ly'6
5�/)�z`�>��;� 7��p�!M\?ŋ�_BO��-Qt�a�BHI�c��*/b�n	�n��V����{��WP����)MK.98]�2N₉�o��!Kؤhq?h>H,,Df��}&��I�,IB�η$d�z$��.L�V�5qa�|�X3��^���q��F���1�<Upٓ����T�;����԰�	���~��hZ�R$֧�q���9��)�W�I�pe��l�9�7zh��i�.>0�*p�:��'�@��������F0y`ƸA?��viL�F�Y9�TՏ�����_`w���|���aυ��[�f���$���S67Z7T;��Wb�.>��u�>H��O8��Fa^��`�<z�Qb����������I �߈�\��<�$�3<�d~��(��j9:�-�k�� ��S/��Q�Լߟr.?/�gB{ �~�5��{�S�lb��]�W�}�����h"zO��1
��2m%Wk�YʯO���ʝ�A�RW;Ӏ B��ó����媃�l��_T�Vx�t��'13���b.�oUf���h�w�[*��ǉ	!-�`ύ<f�T�MXʯ9�3+T+�t��=ƿt�K�9� BQS�η%�����l�@q�)�i���6 ��	�Jʃ�gF��@	N���q[RN�`-���_�0�}/�Q�TK�5���|V�l��a�p���w�c��7����~[c������Kv~lƮ����o	~��B��O�ž��/��췞�-���Z1�9{Y�Eq�^*��M��=	���u��N��V�]u�3�8t�<$ǝB��eD�7�C}��f�/�4 �yx�c13C�,�7uUl���20�=�A��8{�F[׬i(��K��{��]L ԓ#u��>az�-�>{���f�������e&���ۣ�K"�����v��w(�R\��4��������&�o|֧�*7"ƛ.�v�����xg�Śr��h�;:ʙ�C���j�q:�x`4��o�� P_t>����*-�<���C��߫��F�+d3W�2��2*lǘ�`�R8���tWrEq#�j����D���'�������^;~��8���<A;HE~d0�a�O�J���v��3Ӱ9>�������w FǮ'�3����K8�a��	���ԗ�̲?r�ix냋�G��e��B���b7uhǒ8VN�8e {��~���P���u^�ڶǸ�C�f^���$Hy��ޫ����h>����/�x�1��E��r:�S�� ���
�ể����5��^ع
�]��������� �:�IuB��k��e7��)�Y���f��s4��J�`�7����丹axɚ�E�w#�d�`j�c]�I�β`�^.����f�揯	�4\�y��|�|n��;����W�Vn޷��*Q�y�\�\Y��y�7���Α���<Ɋ8�:#Wm0v@�<_O\dDu?+��JA��s?�F�-�n��}�R�R��s�� �8��������zz��s�� ��2W�ݑ����C���҄���pг7 �q�n�A?�2�-g=��N7d7�s��[�rY�3�ؾ�9�ud������iՕ�?� \.nPLVG̞3?qv�?�p|�7� Dv��#KE�ꆍC9ě5�$jDW����.e!���[QM ͈�}��p4JHE�xʇ��Ts�?�I��q��@�-�}�f�}��i���Ңpf�q�����`^z�� e\˖k��R�L�O�8�ff������F�}�_�0b�7,��Ip�����b=C�����H�#O�Q��-��ư��kLoo/���ە��s{�b�~�a��J���A�=��<[� ��;q$��n�@����=��?BC5����$f��QD���i��x��0P�S�/ZjT�<k�@��J�aJ��ЮJ�u���8[)�I���|��~��G���e%���w�(�������t_2|�e���ȫ�nC� ����=f3�4�d�j��v`�'3��7���u]ENi!��āg�W�n��t���Ԭ�i�[�y9oK�v���C�6He�	.�U�^e��:����O��:���N����'�h����v;(k�l'g�gV-��;a~t�n�v�A�q���v6��� �c��7��b����*t�k���߽C�jS2L83[?<��^׋��s�����R�_�/<���uE����♪[ht*]t�yq������us�x=�z���J��wO�u'�U�/Fj���F��RC��C�����ML�(%��]��^"���Yۥ/�~y����!9Dބ���M�Y��|�1�9�:cΤiXly���eb=�T�hԡ���5L7l=f7d��(�c\�/���8 X��/�	��㙨'p��خ7:��*�EIԒ�~�B����x|6y|S\vF~2|]	�E�Nl�}\���j�aw�c��s�zÅ����O�F  j�;6�F��BuFӏ��}`4%%_3
��_\6/%X�S]�i�7N�)�H>�4�}�oO��ؚ��.q��`ed%�xۆc�N�v� I�(�#�
D�d��~�����딽;�>���mG ./_��&�>�2|j���B���`\�����>r�6���,����y��2�OI4��@g��|���h��[�@��+	ƕ�Z�hb~�J�w1���czQHD��w�2o2�a�z�"މ��%ϖ�pEQ�>{n'�N`��ax2a�:��,$�D��Ϣ�6#�(V)n�����w�n�q;������)]��#��KU�j��F��'�&灱��d6��]Rn��=����v{Ӏ�P�'�u�W���FH6�G�LEEO�nM���v$SN�]��L�(p+#!�]��KT��3@�����_�"ݼj�noX����ь{�Z#UI�5V�5��|��s獴(ڍ9	��(K��$� �����7��SE ��a������櫯����4�,+^F�j;~��g5�5u4�e�A����{���c���Λ����A�n|�/%���W�j�|� V����ֵTCd��j ]��d�$�Xh�l70_ޠ�be�Zx`�7�-;p��@ 4��%��"�x�+�)���ˆ+Z���k��/ewY�MK"�����X)�����ZY��ʮ����9N9�6���W�!Ov�kN�6R-)�E�;��T�Oj�k)*���RCf�j���8=�'�G�e�f��C֑��d9�ِi��H/�<���e�~�e�t��L��.�^�\!�U�&��4[4Ԗ��.o�֝��(`f�a���9��+�>: ����n��US'���������S�=|Җ�<=���qč�[WA�l�`6�CL�bb�$Y{n���^�
;�WW�@J`�|�{�1��Q-T�ҢȣcsQ�9��^�&�oƹ�h�4N{3�������:�1ZP�'��庰�V���������.�u���`��.��n
29k��X�jV�Imȵ���b,���7J�P0jx���T�'�;rvvV���\��a������.;���7	��O,.xSR�ҷ��J�s�13�洴��j�|���f�������xPS[�F�xH�� �F���iXi�=���<_�lRH��
�ǃ�r����0�BǊF��}�ݠ�겹POtP'�<5�j:��ZČ����_��
��''+��!����EG�?G���@���VRen5��D��d��Z B�Uu�ԗ5�$��MP6Z���`�T�ti~�P�3�iSTz	������v2��2���m����O�pҸ��U3e��[�Xd�	���̐�塏���������`߯��O�-�:�R��c���2�A+��@��ʗ��4�߱�GG5��I>�D�en�L�aǡ���ϰ��^u�i��	�_���p� �GD�V��.�s7�.� E	5�e��rP�Y��i�^{�5%�6�׿I�_uf�lH(j3�w�'�̽jAa��_ꥦs�F&̧�T� \4�0��|����դ�s;�!���t:e&���ԝ��^�#�7�<8٭��Z��E�ּ��0��� D�@1/�n�ҟpp0�W�0@���F���֩ѥ46ukaI�q#� ��(�4c�}W����Ia���/�`�/~")���	]UI'q�a���r���?$��p{�o�6,B�_�ك��.d�]A�W>��}�t��`��ƃŧ���+����r�/Q�7ׯD�x�J��O(q}��&h	:����u��ݱ�����r�<Q���{�o`c��?L��'�H�
�RG�����	��y�6<臍����x�so��H��3��"����1�� ���Ζ��Yn�l\Ȇ�����.�rd
1g˴f�d�3^l�"LS��O�;Ӛ����P^�x4Ʃ�$j��ߚ�XG�q�WҬ푥‥U�4P��jĢ i/9%&[Hsd����<a`3�Y�bg���4���x9��n��4��BK%[�!K��_W��ά*�#��x'j����]H�Q�]��Ϋ?yꖃ��Tu[a� �"�!h���!�D�cO�瓁�O��丒.�Y�bdB�!�����LW��~ܐx���7@S�f��E N��(����.�s�"X�'�O �e�'>�챦�D�6�q6��G*�$��ta�����Q�*9�tt��֊	���xd3���fJ�Ї}��"�f�vPy�r�&351��� /3@˓8L�h2WVW ������4�ͷ}�>k���;Ϥe��`� :��:������̎�����i�<�[����	{�=����X�3������1Z�,ե����m�(�o�M��ls\�|3�jL��%��L,l��+���}��S�䰿6���B+B-w���)��ڼ�S9�u�_�[�e/������Y�:���,Z���n�!�p�n�8�`����vu˨���\i�����?���+:.�y����<�e�@1�Bݱ�zU�\����?��W�M�����{��~�w2�3o\��	�q?����b��u~fٕb� x�v7M��Ɇ��V��H�1O�s03�o�:đ�af�b!����x�ת����o|;�k,0��I�w׭�3A���.�� 
!*�fۓy���Ǻ 
�jd� ߆�XQ��=ο��4Ó��_*'�f&��7
v2ƽ�K��j��q���ޡ;2�������v�� 9�6<�E+=���yPK+��+�A�f)��A�����>�kjc����7���� ��`HB�]r
Rl��������%}V�lUm�m�G���k��؆�~�E=�h��P����֔���e��k���^���=C�yf�6�����ݎ(���s�<�Mآ�*�+Z?E�g n"�))�ӱ�ڍ`�O፧[$��Q�GNh�������7��SǕ��6T�@0�La���.���j@�
�-��,��`bu+�o:�Ə=%��m�-x�#�_gKN����e2�e�{�m{���E�#j���/��"�d��,NF
<��e�^�s���©5�Y7w
%?y3�+1v�#��Ҡ�2�o��y��q��"n��Ei
v<�0�_��DvbY)g8�m�E;�ʌ5�����N����#b���]j �������ހY*���&����$��+�w3��^�j���_i3�=O\��Z
�Wk�b;/Y�j��4�����Cn	�A{<�Mvu����q_�2���I{mZ�{����'o�jhא�����d�EE�F��~�gfA-�`�]��������B9^����F(�mhhK�\�]�������H�*�搲��� ң�4̓���={�����_H���bc��Px��5�ZβP+/��s�a���-�j���}o$>r�O�_�������:)�
�)��T��џ���|�5�ݶ�P����H���*3?o"���7o������b=�'h%�p�)#���5��'v�8�3u��HΟ�w��ђ�5Һ�;Ms 8���ʴ8�G�
�;*�[�v��HS�~W�ʚH>�~?X�yct^����m�RP1�"����䁌�����B!Á�Z�F�/ѿ��-�初W+y��[:�J��**g��s>�aQ*Q�����tn.d�΁�����,
4��W|�G�E�Ue��ܱ_��EA[
_�e�|�)�/����c�X3��6�=�k��q(|kn<g���a����߇sS_��D���D#�74��`y^�1��X):	ޙ�>�e��U���׀�AL2ָRY����h�v�Da���_6*t�p��cK�o:�Y��ص��*�W���2�1�v�}}�D�[h���%���g!�M��/~1�H(����?J_X�Jl�|�ɣ�ʵ�1!}8�6�x<7��_�r��g������Ss۫�"�sK_��R}����sH�I�����~���%W> ww�F��B?_�E�1�%[� ��k���!��c�?��G��]l�*`J�CC��7"G"-�ܸ����h�ծ���*�r��3��8낂��Rk�ԡ��x��k'��.e+dSg"�O����\�.������@\��`���GI,�HV����Ns�O[�b��`g�������_(�R<�ǌ�c ڮ0Q�Xj�	�
E����w־�DI�f�h���`Ux�g��l���֨�����Cyy@m���9���)��L�����ݕ��#bgK(����[h�ä,��f7��_Af�S����#M���:��]+�6ȼ݁s4w�I<�:ݴ����C��7zw���(�걲������Qc,�^u-��Π��ja���w����}s9���*,M�{�����kz��o�us�4���GyVD7>n�����sݸ�n��Ţ,&�L�N,��RH�.��a`|���D/^��V��KFju��\�O�۠�ƃW�x%�8�b���"k��n��`,�fݿv2�G�:��Z�f��2l���9V���N��3����fL�R;��>�ӚUd_t��&"j=j�t���,5�����0�.0kf����\�Y0U�|S�k5���)[��&gJA:1�@Qʷ�Y��X��$ϩ���#�fG�Ѽ�c�s�z|����R�ߢ+[���gOf��M�� ?�вcG7�[���o�T|�������?/ƤdXҧg��\Y?��Ts�B�3��%�����`
����9 'S�:��|��)�-L^~]?� ʴ���v��c7�Q���U���x-�z�е� IV����>2�#lڮ�fݍ��Y���G��ޖ��l��:;<x�hV��e�%�Os��{��o�X�8l0�� Q���I�ն�)�Ǔ���7Z�e
*�� ��˵Az��~��7�2��Ґ���u�=��v\<�\|��]��$}��Zp�2^��Ihi^2�ȨJ5�P?K���0_xں�B�y�`I���.t�g�
�k9�*�fA�fҪ]]���73v�ti��]D�쟮}5~Kc�4�#�@ߺy�qR/�%�՚.?����n	�ƽ%������L��H���f�p�l0�:4����AL!-gL���3��9�-�¦�;mSb\R��q��L���5�ʿt�hR>3����2+}�b�H9�?��,��m�"]Zz��u��
�z�#Q���`�/�C<^@��95CV.
��WȊ���4��/~���$���~��_�N��U�,"�|+t����p�	��]�eSCe�fB��@*���"��:`}H�4���F�P���Ο���F����:��t���Fh���?-dl#��Ub����8�O�9xƫ\�%Jgn���5���{ɓU*�ö������|�m�_w�R�ɬk��ڟ9�|m��~�iK��&�K�58���}��*��k�[k�kt�C|�M�a�S�<��5!��6�r>�c��7���H�'���ٍ�=�i~唵�w8�Z��.gB���,�aƆg��
��*�< �6�_��� �n�d���[_�C
~��任����aƻ��M�e�(QD���ڴ-����s���>�����Z"�x�~���<k�����DP����#��o���y,X  ?��iN��ݯ�-�R�=��R�J�rI�T�OH$ɜ.6��BE!QE���\p	����Ĭ����,�?6�j6[Ԕ�[����җ��%�/�>iq"v�ܯ(�Q���XH��yx4��+���[��줁q�i:`.���<�2�40#�S=�`�����/��i���V^��v)g�u��@���;9�l&樋�LÓ���{JFo��{a���ٔ�#%�*$��NL��/ݐ�+
<��^|�/�$�xQ�91����!��c>�8�5������Ӭy�C�tABh��Ƚ�ZT�n��xer%�ռM�?v1���Z�9����Ot�6�S�[ڀ(
�wUP+�K�����������㑃 3�^k�Ͱ"t�G?�V�J�M���o��%��##O_�{'�НLv]�i��^�3�ۼExq��M|����7P�	���2�K�4�.��z�x]6�7=rg����5�nE�к�y���Uvd�pyP��bC�1₨�ϩ�!'�-�fC���ɓ���Z��I�2Rj�h*.�AI�m���ZWMM����e_犰`�̕2�cq��Ժ�����(<2 Q������ID�R�����TO� �-2ۨ�ȟ��nZ�֞���2�*�\��ÜG��e�A�x��M�c��N}���c�-�6C��x�*twS�Jc9!���Z�1�1�/\�t���-Ul	�!3�8���t��BJ���Ҡ���d��{۷�l4===��T��Nm���'�Hx$"!0�4��qm���������s�kT�0���ָOt��Kf�e�X�s�(��"o�,)d�����襀p�V���r��n���ٷ#�rK�O�=�#��H��
��Dc=��A���f���19&8��k��9��i		7�Ύ^un�]��^U�=����p������ʍƅ�r�U��~�m�oQ��8��V��F�7��8���D��j4�#$�{^o=:E`�3����7�����А��T�>P�
i)6UT��k��+�j�p��]����k�3�V���sWY���Y@A��e�̋=|z5����AS���%�S�z?1&��?�6`��1ǯ+ G��S��&��-QM�*
2b+"�_Ⱦ���<:n~����b8q�9���bW*��+/����j?��|�J�id+�-8 ��-��K���JUH���[D�(.�E�j�mb�V͉Lc�Lh�u�y���F�TQ�G5�t%���Vtڬε�<����s�p5\<�zv�SA NQA.dx����~'�֮�kh`�d(J��Р�x�23��v��58�bF��X������r�}iaP)�#��3�l8�IVGa��S ����dR+"����x�&�*p�m��5�����|G6�;^6��01ԳXle�n"�p��	k��,�r�n.���]L�2x��<<��<��m|����|�����_�*f��w��f4���*��i�s�o�<4����4�LG��PZŷ�m�9_B�G�%NU�I��@���3�����(!L��\�e�����+�&%'��g�A6�>���˺�n�a�8�����Obl�~@s�*���ՌGaiõ�j�c>�q�,	+�\�q	�:={E��Q�G(5(v5]%Rͯ��P>:��0v�/w�e��#�~Ǳ�&ͪ10+�8Ɔ���uC*e"{�f��ӣ��5D/˝�s��p���o���U��j3[�fHj�LA)���3G�4������ln2ۀl;T�u����GA�U�&�S���Hڣ)�p	5���ŝn�H���J��I�''%i�#-D\N��������GdK?s�T@<2�e$
������-:z��4t��a����U��~ѥ��J�Z��c��%A��HG���B��&Ria����� �%�.3�zDgub�?eZ�`TŔ��O��sF�41�.NF���s���%O��9���0�a�۪B5�Jee�č��V.�H4\=��[(k� ����f"��n�+���4���v��r7������q���R������7$��}��l���#�ü�
)�������Q��<֘�$�<֩��2��Ȑ�{ꭵ��%������ykR�8{�2��>\�C�:C��(~���)�U@Zd�ظ��0��dx|�����Q��9T��*���Uk�z�v�+�B]�y�AK
B-NN�&Q�4�L���ܻ��i���VE�]DN���E�iۆt�`�f�>�qe(5&�Iݙ	u�켱<7&�) i�q?�{G����?w��p�9�0��C8p���W�B��������� #j�*i1�~bфz���U���c�W�pFMy0cr�z��ڥ�'l�����G�Ƭ��/�(9h��Uo�]����U��4�� !r�=�#����M��`Ó9�%�/�N�0\l��@�ae}��F��C�e��l7�SPR&ϟ��z�-8�O��H��d$ͨ>$��:�ƽ��Eeȸ���>l{�[��ǴȮw�RFH�<'s�9WS*<��_y��鏂��ą2��E�����s�C}� �	a�q���[m�;�QUK���?g�_&F��Iܞ��X�02�\���"�H��b:m1�㟃��k U�ܴ��'���_O]τ�A �J/�tA֎�Θr�|�n��G_TCK�7%2
#O�gOKZ,����y���4"NA��^["حf��G���yU_���jJ�� ��P
�Yejʊ��+ZKJp#[w��mQ~uz��ڊ|�ʲ4��L;�9� `����be�
A�?��l��b��5S�D�壯.x]�an�kĆ���"��T��P���zvd��G�#jK��yR�s��ݕ��� ��b�9�v���׼�u����I9QA�#5g&1 �л�-V1�</=��9���N���&����AkӓC��m��r�'? �}��n��ǀ���RW��欠C�|�k�y�k$, ���>l͉<O*�3K|J�Q��� \#����]���#B�|V���7���3�~���=(Q"�c�n�ǓwM�\;	�o��o{jk�bV����</M�ae�Ck9E�R��A��Du�B{�Ƌ�=��~%6�}Q�5��b�8T���J�5Bt������8�4�fK���E��0q^`x��w�D�ۗϗRY�dO`xм_	I��z>&S�,�Q��x�͒�W�/Ip����Z{�߿J�zjx��G4u_�!%���`�JW��i5�d��4jC��I�~���#%"�Y{���V�,fq����)y �`�Ƹ�`Νh[����IO��T���(Ū썍���&�4��n<$g�G�sd���*/jpF�&WJ}�R�����Jv�1�3�dK͖�,����<o�I�I��S_��6R����?z�{^�޽�C��^��ԝ??�}�y��m����xݟ93��Hybɑ$1%YJ�����#���XF �L@HaL�ȡ��#����D��n��׾o��=?�=O_��6�{����/�n����wQ�=���9x��6�x~Y��b&���N��I��p��w���m�{[p��y�}3&z��p[T�|�[�P�Ye/���x�媦%��!��X�Ӵ�@&���D۵�U`^�9���\I����ht+5�-fǕ���/.vn���qN��t�IVT��0�f8�Ѓr�f��w�����$!�M���������HW�4fc��,��c��ki�������e�}&>q ���u�&ϽA�3�djmc���nq�k��N�!)T�_E�V�*�/Лpͣ	_v�1�/�]�(�0m)���?n+��R�%x��E ��{D���j������ �(STg�Pb�s����=���,�tL�N;b@< �e�����).	��`��:��Buf�j9�m��p��i��g8�pu�9_Ǜ�7�0��h�3�WT�/
�H^4�����Hk�%8���������/q�/Q�q�5puw�b�a�4��K\NN�Y4��`s���m�ڴpGdD���Ã��f���]o�ϓc����{��Ȇ����-x���_w}	�j|A!^�px��){Ln@bVq||X��Y��̑�Z�9�;�����WHP�tO3f�2U�FS��jd @ˤ�����j�J���"�_=�t��^����:��2�ʍ�9��HZ�Fxyv��t��W���മCM��P�C��x;je����HD �yI�M�h5l�*6k���!e�FS=d����4�-���������,62�$9;�ܑ�׎'�u��� � S��V�U���x;�3����F�Bg[{bKLH�d�I�}M���:}�v<�;���n�{ٜ�峁�7� jRPT���< �G�a#ʈ��x��ԓ��;��U��fP?�,���a�����ndi�̸�8}��T���0�������)�~>iz7dv���5��髑���?J�	_J5=�\PDr.KʲÖS^����=.�"���������,7���o<���8K��I1�.?���.�`�Ľ��Rl��"g6��v�W>Ĺ�,aI}Yjw *��J�[����?�9�7P)uz�dQTqv�!�|0�S���xԤ���ӑJv7O
��%�D��4��{�}T'�Pb�2f�]Jj���a�vfyԮ�ȷ�����F����Y�P�q��m��c�Ŗ�e�L�O)�$ɔ��e��p�,����>�DS����� ��ȊZGz�3s�x��k�Z�2�2�IS�h�E�o`����2{ s2��t�,����[K�2ȳ�-G�nb� �Ks�6*NZ�4��ĥ�*��;��)z��92�+��E��ۑ����/{���9<š;�s���v��P���f[�%K�P��֟IuS�d\h�^��	��UݨQޤܬ�Y�o�ݗ��Cox��6V���	#�c1M]\T@=�ka�Nb8�=�f�h"Ǹ��r�\ʮ�_!�q��]h'�5i:�Է4 ȓH�`i6`g\�y]pS��*G^Ӑ3iT��{��2q(���a�}?�{�ܠ�@*�k��g\��H���]yn���8:r��ڀp��ZX�9�����ץp�٢z�A�GZ[J'+�����k������3���lW%��,����E[�����#�c[Z�9߲w��`�(r	ZZD~���u�Zf�V��<�������~+vDk��֐�A��ƀ�u�-����1Gs�#q�Nd�Llq�m�1�N5��t�z��"�^�z�9@���hu7�nL*/;S���i�I�M�m�A+{�\��Y�	����YzL�f	�5�㶟c����`�O�g%~�n�K�`,YmDi�]x`�E]2?nA���8@������[ΰ��£�*WQ	!jw�D��kDC.�L��@2��͝V4U�c������g��RR���J=�UB�m��/�U�( ��~��^t�N��]�Yh;k��^�,�nU8n�=�F�nE�X�'@��|����������CƋy���(ܕ<>�@PvH'/�i�J�&U��0R�=^��`�HH(����*b���k��j�()�����l��̅�EE?����p����`���ie�	�:��H�w �g�A4e���?�3|Z��ˢ#TtoAPᖥ�� O��j�`��@PZ�1�۫3��n������.l��>߆��\�}�,���k��+(;>������<l��oS���3�9L(��E"h6x"���[����(b��һ#,	�x�h�H\lR���!���|���}K�L2�D(�"�zD�l�ݗ�5�'x�.��a����j;����5�ʙ�f��Q�Z\�~�������^p�,tq0Y�6e�s��b�t�5�H��p����7�j��c\��>g���U�u����$�3a.[�m��R�?jPr��J7����X�(
�i�	.B��%��)�e'���@(3��L��|��9�C�Y#U�R$���P�dķ:��[��
fg�J���8��I�7v�����h�u��7�������A;_�̙�ñ�;��}�b�Z�����,�%��Ǚ*K�����K�n�5$�������ݗ���W���E���2u���`��t�@ґz�c�!qD��Z�d�Zq�B5pF��	�d�z�d�5w�}�!���Q�B�_b��տjS�;C�0"�}��6!\�"����t c�4xt��EjB���m���M�f~�sg.nE���O�赞u�PF�kU�l=�2�͉�R�'�o@]jk:k��*g�!��Nljz�Y��H��M�ΐ�8ɗA�%�T��?j��`�dTx��i�gi�	��}.�2����H�	��Ue5u�O��4%��al4S���o�L�m�i���2v#)گ'�����"d�U�P	$Ȍ�6#"f���V�Y�����{�wK%�����C���NēT���'1���۾�I/�#��:[��$ۢ�l�w�a�)�}n��1�c�=Q�{��,i�/n��0g��I�P�,hM�ҭ&ف����C�D�2�}��}%=z@���UW���6�1��N$\���i`�B ���<�����?~����؈=䌝]K���З'��@�!�X&>yl��T����aYk���@ى�t;��49:E�k�C̟�Z�梠�h��.����x�5���W�_�A7�ܺ{h������v�,QI����*p6�&�Ă���l��i�hJ��PŚ%�!EQ��2��E�F���*�j�[��ޓ�e��4�S ������8P8^�M�;B���u�G��B�Ngm�Jk��#��3��o�����s=�M��B��/�Ne����⬵���KD�����)$b]'���	RX}ST��2��*Ȟ�&E�)�E��J�A_<Ït	5,ۦ�^X?��F&����Ir�Jn�Qu2�]Y� R>��9مo���B<�|�& wAx+����\���ClM4
'�������}�1����Q?"�eqw�>�k�^�ֲ��������x߂n�d������GZ�,��5��Ϯ{�ȳ�tc^��=�V�i��Hy�%���'2Ǥ���J�T~�u�.S���Kn�MBC���k�I�`��kRT�Yp�xid���8�KJfJX��ˤ<L�Ta�wr\�WpQukjv��Y��Q��8�M�N��|���3�,f!W�x8���|�>�N�<~M����`�-D���W���#�<��Ǫ�.t�sO�Ѽ��1�g.��A�JU���������݀�Y<K����оxǯ�#m
*o�����3�d��l3�^k�Ϻ���k�!��πp��/a&����i�N��>�R���^;��j�
�$>PՂ1��N�J�I���M�@�7y�p�̪�
J֙�*�+��e�'*��F�@�{���p}븟e�QD��q�������y8�:?8Iɀ)�.֠���,�� Em��{,ML�鋷�lY�܁lm��ܗ�_�s��_�K�с�UO�nXq$��T�2�QU3���9"B3�RAFBd����7�������
l���_o�V�m�	�T��
��1�<cӧ�؂�Fj ��Q�V��d@Ƿ�����9Է
�uB)U�1�����Z���l��ڢ,��\�3>$Z�@��mT;���������%�u���ű�%��%� /i("�_����ׯ=�t�U|b���~ �J��i��L_Mr�M�-�Q��#rD���*�˚��ld�i݊����X�����6���z���h[7v�۶m۶m�F3�]�U���1c�9k��}��4�@�������$�p�$�����q<S�H�Q�ƪ��)8�kY������q�����������C<44�����Qg����\{NX�$�G��-�Qo�:n�;�6��e�w!��EǙ�S���5"����L@ L0�V^1�&����{���35cXPP'{N(rOx9�
(h$KzT�r����s����#B�Ҹ�t�}�z�˶9ĩ�Ҕ�����W�a� �H���ް� ,�u��N�E.�S�Eu�+s��V��_�C�ܡ��ѷ���,�t�?c��{��H��� Xhx����Wd��Ɋ)�i�\�����ɵ��˴��q��9Q]�m�U�f3�2���-�4��X�lc���C��y�M�WAJ�	��OT�r^�L�w���P3w�w��R�<�rs{(n�D�{ţpA���>��)n����O�E���H��ʠ���^V������ز���ƺ]"���=AN��i�ο
�T���E��RW�'��il5��}�s �25�{����	%�}b�fSݎ�$׍m*�Ŵ
Ƚ��f�QR����,��ߵ(��|�VH�l9Ɇ�
F�5���YD���ce����9�I��u��3���8K@C4�P]��n�f����g��Xe� ��Cg?����s.R�c���H��l�R�����Bp��	��]	�K��8��Pw~2%��6<��+!�/仨Zl!)'�1E��"��7��To�L~)�E�l��v�X���kO��ӁE�ZQI:�z�¡����2թ�F�4+i�#���.ݝl9��� r��茼bԄ�vB���Z����C1ă���냳��)0ҿ5ܭ��UV��'+���,��LM�t����|ݾ���c&5��ɮ�q��'u��7����ȟŅ`���֐&#�&�_�Eu�	�R�-�l�e�,*�͔���nˁ*�sH ��M��Yp���ǏT�d���-^�[J���!�X2�4�Swߺ$̈́��6*K\O��Ug��.ί���c0&�c���2�������'9�ԑ�8�6��dr4���@�����ǜ�D�%
.4�)�n�B�Li�E�踐��k�?�W�|��~�dXs�M��U�_�r��~^_X���p����=�z�k����"8׀����Ʊ��n�}v@����[��2	�s� g�K,�����M����n]�®�Т�+���>-	��F�M;g���C��$Mt}} )�����*��9� Q�QFQ1����_���ě
��˵�P��تHCN�w��.�"R˒��[����J�/�"��X�o��_� _a�,=�[U98K���Yt�֤N�Z���4�eQ�8caeG����%_�G��Մ�"��+��,y��f�SS���(��q)�SC1���C1���O�F�4�r����z~Ӗ�����f��vBw`3.�iƐ��j%w��un�f�N���S�ǐ*E��H�,U�u&=�	A���ߙ��z�	X"8۲I��y�H�����=Ә�T?-0��J�iR^����VM�Q���L9�W��)
�c�V~��QVY�X&f�����k7t����YA���Q݌x�S9NT�k�����3���mW'D����=����˧F�ŀɂ�\j>l�x_ׁ%x݉���=�Y�IPAR�������+6>���)��mznȝ���;}���Rm	��AI/H.�'�o<�q��r��UAB���"$��r��|�J��_�M�IC��ka�k��li�wI���j;��F#�k�0�j�*�<����f�q� ��}'��ʒ��Ϗ�$���zc��E��RR*H�����&�zE�&X��oX��eܷW�X�~̂�fC�Nk����<�
�;�ɽt�=S@�^��{���t'9��]��ȩ9(K�����`��V�l	P�DqN�V(�e��s���**x�B�G���d��5^^"h}�v"��4A�HE"|�}q�P�P�#U�U�^.�H�'��Dq9m�e<�9S����ߚ�*:Ջ�FJ���7/| C��H�1��F�g��ZS��CMI7��ٍ߹{϶�[�z��~t��q�T�n��/|��7�*ˑ��ʦ*ׇ�)˖�"M�ce������l� ��r�폴#�;
I@�}�mλp�8�R�t���"ۆ0�����t*��%sq����ymz{);B�����u��ix�������@���G�~�b�tMΙ?���[~�U9&�;�y�)�~F��hk�& }gҬ�D��N��+G�^a�|ح.�����I�����	��&)�L��p��V��PC���.N��P����+�%[n�]�O��#x�/���qtl�`�����9 "W��T�C/�E�C�x���V���Jv��S%�'��c��+"��yc�pS�>¼���C^{!���$����[�Eyq�3q�Y�$߾��'Q	c0Z�c�nfN�SRiY�E���i�X��
³�)#AJ��#�h�����,�H�4����}~�����'��d��:�M�l`�+*1jC�K�%|����~e[Q��`���ߪ4���}+���~�w+�?O\d��w��p������HC��gGq}� $�{�uֺ˚P��a�D�������:���;�|]ߑ�<� �_�z��U#�mb�z$�f�&�v�R���j��J��M�%��ȱ�6���R
f갡�dZ���وP�������!^�X��e������]�6y�b��5X`!��k��5xv�%��.���%[,����sb�>�@V��C_�����OD�@��܃3���l��Z�C^v+�vzG���ڄ~)�����7H��vu��D�͛��5�~L0sB���V�j�_��c���v���Gq�F��]VHB���X�X�#K���f�Ff7��CD����Q�A��P�IE�!M����`�2(��n13hLY�J����n8 �Ą���3���*:#{/$�̛��i:�a�޹[�G��^w՘�`�TFo
�U׵��p
�F����q���#/l��:4H�����ug�>��w�	��jkF����	a0 ���O��v	p�GO�8�����?�J�=P.r#3c1\�����6�D�}+gնī�S["�B��z�?�n�۳�}��y��B��AJ���"hvf�f��&�p���kz�h�u?��(h��穔�_��b>�؊T׻�QJ�g�?u֩���Is��f��з�}Q>�`�h���mЁ�'�<x��`��4�H)���z���3��M�����x���-
����|��P���,�eMY�j� MOQ�(cY��q�'eC�m�h,*�-��NRC7�����AQbR8;��:6{n�[`�lg�PL���Pu��u���L�!�#�<v����=����R9N	�?W�H!�#��R
��We���QJ!k ; ��Oߓ��9�eaF�:PPf���T^*{:����#^«�U���� O�2/D+�4�<�7����|�,y�.�;���q��ːOK�����QO��Ny��	��@Z�0��
�Mh�x@�#PI�[���i��"2��d�U�̤�J0��a�����beI��NKlTM����"��4���(Lښ[��GgJ����L!��k�Ti����	Lڌ�o/tX�A"�@Ā^���K�&�F����Xz)б>,+WΙ���Ң����K��6l+���f�&؃�m�v�$�o읻c���(�g-ڽ:S�6y�����-�J.ĤM��j��3��#�N	q<@�W}F��n��`�	p@��M������LS6�I�T($EP�z��c�Z9�޼d��v�ֆClҠ*W)/b��af����q��xH6�`m���e����n��0�4��f�}��&#�>jy/�9��Hoώߛ8ʪ갠���O/>�6� �^��sϣ�Xl����#�E�Y�;�]�)wE?q�����}�Ԫ���Ҩl<���T��{=�-��Љ�V�X(��>���~��+����*�TKJݒ��W��#�_.�X�c딌E�4BU`�.��-��$9��xg�Nw�6?B;ifF2w�Gx%�|�Һ�*���S���*i�Q�aX~�����-���O(-�+(ի�+�'�J�=<�8��Äh����̪.��}<L�Ӹ���y��O���)3��>���̻#��&�"�U�1K��O��E� �ʍVIo1�v�c�lmD�=��EA�=!�/z��F�J��炇W]u�^dw�zm��tK���K�˚$�h��O�&�,����ٱ�TB��,�d�܋SGş齏����>���J���*5;�o�˰y��?^B���
+��tڏ!�r�zȺ���E�Q�%�E�0G�_�`2�%	�j�X���p<G��=؜Vh;V����݃%�ܦ�m4�i_Ei8�Z5�%���a�lV%KVE��rlBP=ꩈ�CkVM���R�VrA*�Y��7tZ�F�΋jG�9,ar!x��0L�ͅP 7~"p��B��Q)]Mfa~y�P���89Xd)eɐ�22����?y����g9"ƪ4e�r�M���h�3��d��@��L ���DD��|��뛔4i�?�2!�p��D���)�@iH��7���9�+��PZtC�m����=�CUse@z��b8���j���{���CC�NW��O�!�-��h?Ƈ��hhȐeX�#������ 3� �Zs�,#QV_���p�� �����֊Аi����ʑ�%	�>I�]醺~�c��7?�����跆>�[򄕧��ә�d8��&������A�=d\���\�"��v!��g�Aآ"/�F[���Ț�����W%��L�Yc?7�Q�6�IC:x����~�g�wܧ"K"�@�J����[|��v��[h~ ��|����&�C��cJeTJ��҅* }���E��G!�FQ~�@��F7˺�j�%��ƠV�cnX.��j&�;��H�����-ax���S��b��6�P�W!��Kn_�%�[�� �e5T��$�f{^2M|��s��eu�\:p.����.'.�8���K�؛,~�m�Ds�������8hn޸0��j�?m��=����� ��^��&���4V�f�6i���&�R ZW��>D�vv>��3�b�A���*xs�(�9oA��r���(��]��Β
��[����K&���n���.
�n\�\�y�P$�<x��~<�-�����x�i����P�odT�I�t-TU�0�2O?�|�~�U�/ "8���݃�g{\\�vE��_:���[�����������_��1���6ρ��z��� !@���(���,J�f��P0�>ʚ@V8��,��ډ�ػ6d�$sγN��Ώܹ�	
E���Ƣ)��mM��#o�����h1N�aMjd w������_�I�C�����i����#�D��C#�!,�ca���2��VL��<A�r�� ?o��h%em��$���$3'=i�UU���x�Ǔ�[E2��Xxu�"�Ӓbf�
>@����hʛ�w��ES��01�ڔ��-�W!�t���9&����A��d�=���CB�I[L���j�	���~����fu�?�y��hսk��`�C��X���t�@�m�-�k�V���g�D������LzI�a`'�V�=��y~E�k�^�3w[�L�L��T`%���7_J�ǇB 8��x;U�ϊ�Y�
�1e��l�է9�%GA>��4�q"%���
I��VŎ����/ԣL��4j�WY}FP�
F_L=X�ٌ�^c撱�lKj�۱"���ԯ���A@�,K������JM���8���t��?]�����o�w��'���e�cŖ(w��� ���b�R�1@ȎO�v�+8�J�N\�.%+��s�\�
��	]»��	Y���eQ��E���5-Q�O�N��f��y�����~���3a���!5��%(��΄�GA�|�ሐ3�U������+ x��u�P�l���a�,a'1�%��q$Z؂�y[����� e�j���]h�ǭÊ{n"�j@��xsɘ����&��)�{1%t���*c���e�`t����\�@��CA�-��~��\/�S���8vFU8\��
��A�S�fܡFC�5o�Wf��f�^�@=��F���ȸ��6�]��ĝ�dO�<p}������Y��h)`�^ʛ�0��>�c��M�j��U�3P��p�<�A�!���^y�n-��/s�oN�s����C��;�F��>�(w��.�7��4�f�#��>|f�,�x^���iُr�~Р=�c9GN
�P
�o�J0���
����+�����(�u��N
{�JF����l��0^�FV�y"������[���1֮�$�K�Q̚'����`�[=@��p�չ�T�J[�U��=C�����VC��G��A����9�#,�5��Gw�R��l�6���N�iP�V�d�KC�V�c�9��~�ydi:�9�(�(�|˦4*��k>}|��+<g���o\�)�]#7�9��^u�oj����A��M����G]v�V��+���ǵ4���o�N~�`�`�rq��T�'��Jͯ\�6@)E�N�ʰ
\��ݛ]φ�.��ܩ������^Y�@鐁R���
�ET����WDL5?Dv��I����S���V�K�L!R���>Z��G$*�;�^����F��7i��lE����f/6�iKƤ������t��OsIqPនF�sј{�J&�G�.͵r�r���͍�-@S7���Ŏ7(~ ����� )"�g�#��a3���_�e�� s���j��"�Ö�F@�*N��7���h���f�Wl�396Æ���s�&o���S�jve*5 �
���³��-QKz��Kv���z|���	^M���X�OHU�=��$H��zj4ع�a
x�64^,��R�{��*���|���������G�:}����i
ʭp|�'~���<��ϟsQ�Y���+4)q
��&��yz����Lyy[�+�l;"�����7)��U�UF]����<:��b^�w�,'�b\
1�-�K���gL(�e��\X�K@�C�e�K��Ͼ���r}���!�rh���xﯤ-qV�V>�Y�w6�*�uf����c��v*��������Wg�ݬ�,�8�������	�������Ć�6�xr��ϣ���њl�0D���8�Սh��Iʞ�1�k�b�+�@v�����n�3FcUB|��R�����d�̊5�	�UNL����&8?D�ߧ�_�1�b�2L�ݤ�m�]т�/"�(�N��;�b��m~�d����	�@�
Q�LXBf{mr,v�_�s�+��K�g�fX�j���������uPxo�6@�o���4�ɝ�6�6�F�[��<�h�'���Re�	O�)iq�s�y�5��G/%\�ّS9���; �#?���`eXV�9sǚ~��
�������#��m��s6�؏]��b�YP_�D�p
x�~�|hI+�u���4�b��ߞA#����њ����m�]n���q�>S���h�P�����7x�7=��I"�O\����(j`�il%����:�,f�U�>8:�yAlp:
�����E-�G@t����� �hv�QR�>]s�{;,�����S�5�g��eֳ�.�࿿*�W��(�c�VR�XEa\��fG��!+��uAT�p!S�����}p��m)�]��9]�K�7�u7ACK��F+�c�BA��K�4�xnNMUXD�T�i��i��J/P�>rϋ��Q�#K�[�OA���7}�Q��᨝>,�*j���a]�!���<g򭟑��w�����A��d]�u���,�/ �����le��}�bάd~����6ڬ��l�㙨�E䳴E
[s�f�!����c��o���y�662��~S:��Z!���9
�D<��,�QBk�b$��n�e
H���G9�#5�6'�N��J�)Rr�T�29�P.3�n.#��\�?��Z,/Ggv��*��@��YO�2j����~ߑ�=������¾>B����mܙ��S~�H}�Y��`~Q�κ<�+n�zUnq!���R�dUk����Փ'����Y.��J���� �X �-��2��M,_WY��"����u�1���:�3���ؚB�V3IN��gD� O���K�mx;#�>�8
�4�U8�2B⏃�ń?��o�?Hg���n�d��t���b��΢�V�!$���ց����^��e��y03�Г�����J�$�s�����WF�oM]��0��?@�a��5��aY�:{�kײ�D����n�Ll>B�(ކ���I}EuK�T�dQ���,L��ܪ��w%�P4V�� �Y4�a��@�"�ZjC��!���~���j��g
�[%B�i�B��*�3�~f�n�����LN��Oݜ67�Ä�$�T�4徶��3q�˽�����DK��)�rmQ���T??��֟�_Xgxw��%SU�*���3��hc��?�����Q�o�B�� �\�#"ժ4R�&����<�Əo;e�lZd�ME&�S]�� D�3}��R������gɹgC
;t��[��ƦG�u�qY:�$�n�,���"��N�=�t��z"z~ۨM BXdk�%Ұ��z��wgxc�� ���"��LDV����$�h��5d���|�����ɾ-�K��}��J�"�c@��8%"�^����?~»��10S��j��&5m,<ٽ�@�:/���G��2:�!��-�ג������|yͣƄ�����O8�UBI�>I�v��=�Ě� ���qT���$��������s��>_d�Ͻk)2�"��P�Z�_��`Gp�Pd�찣������ʂ"@�r�&�-,x�Îr��j#Z0��Qu���6�Q&ڤ3��'иh���m�!�0a�{:��a���@� �p��R�Ί��!ZT#���Lw��YX͛��j]-_�"�䄊�R#O�`��Y�:�-�:y�H*d^"Tq���h��(+@ʰ*��]R�$�4t���>	�f�`72�$��F&�%�J���U��x<�0K��.,��_9���S�<eKC��C��z�W	P�}�~���c�[^B�
�5����/$�W/H�:ɼ��T!�uu�D��we�4���D�5�Mo?Nɕ�*��R�MQ�p-�C9*+��j�^�ph�lQmv�HfJ��j��o��ݐ$N��&t0ښ��d��h�S� �ӪUD�)��#���x�v��*]Uz��e��U7��V#n4�#wI=v�2ȼ0h�Z�=�p���}�&�Ϙ:?�{��F	QcӳB	��Ӳ�mJ��0>~�<�WSY��e�-d�?���'��\n�6�S�Q�{�h?7��Zt#/F6�N컛1�sO/1>��ؤ12VQ��Y�c�S�I�#�}h..j;d\����Т��:c���%�P�����1�����+枑�HkP��# ��i�	�����GI�V��tH��c�-$�����zP<Dȭ��ˑ/����ɲ�Т��1|�),�����6�(:(l1������*�_��o�RKV��du���h����D��'��9��g�جY Վ�"Y׊��߲�b|�%d��e(fX��FT1�)����_�~�:��,/ka!1WW�,~H�����$:A���uj��Ȥ� RͩSM���f���8O;������I�����^�Rf���-Y"�b��w�*�ru��C��E�j��-�D�i��W���YG���l���;-9��&L��k��	���2id��f�>�*k�?��e=���29qq��J��J;�y:po�����P�,�ppkPj>�Q��WA����%��=�T�9=GS�O"�c
�HFՃi�A����3w\��5�c(�p|r{8�;��8��t�A��h����m�N�Nf6��c���E�����<���EJ�6������_&��[�[�����F�<˓Q�'�K�OC�/o�~��r&o�pWl�Â���{x*�p{�sf���49\@⠂R٭�D	�?ڌ���_����3�o%���޻� ��ȃ��:>��<�8ce���7?Xt�Ń^��	����}$�CH4��U^�8=��Bfڒ�Od�<8,G�:^d�L���p� ���M��~9V�����d��O����Q&|��(2O���
XEtss�!q,-C��ȩ�gdF�p��z��*���J��pٌ��aa��r^�����*��7A_�I��DY���E5@=}W��c�U�j~c'4)�f2I^�Zz��z�G������y3��"ݻ���; ����\r	�����^�<_}2,bs��멂>�>��b���.�<���v��R)cdh(�Oz�TTP U5k>;O�Um���#���qi�u�"��xw�����:j��#�c4��lB�ʈ!t�'9��nU̔��<�I�ނr�̋�K�#���p�X2�ٽ2G�m�FK��7��B��z��������;P�5N��P��
�p�ΐf�4�î#���Q~�9n��d��sn�e}!���\Tҝ�!�O�Y��*
��#g�6������$Ee�Ug�`H�6��[��UQ�־o(���A��Y�+��{���Q`�(�RVF��Sj��CK��с�R�ȋP|d�i�x��$�L��БfE$�E�T�7�e@O+ߗ�N�)�5�,I@�5��wwZ�k�����!~��#�=�&�!��8��h�w]�����v�9�:p���[C��`�o�.s��n3����1����A&��}��以r�<���"
nF����:������_I(Q�$f��^%��Y�8�܌w����Ɨ�>J?�i�:ç����=�������N�����!�r���{6dv��k:��>�u�4��x�E:�$�D�Z�^�I������F|�_k0e�� ���Lѡ�t�@��n���8�/ń�4�9���F/��j;�i'��t�ٜRE�{7=������ b����[�w�b
-dP�$�r%�y  �������ݎmq��R�F^)p_Yo2Zw���� �與����5��0�`9K� ��v#Yx�R�m����u�]��O�{����=�ڀ�2��w�z=652�vx%t��G*0��T(P��9* �9�{Ϣk�
��&ըK�S�2�uٟLe(�dE��a,���Z�V+��L7o�芠�>NUM~Zt����vF�F$�&e���*��K�=ț@�q*��u32S�!Lv�n�x�*��ZGƩ��H"[V�/�(��u~x��j����g�W��"�ΰ�WY/�}g�}��*���+���}h �d�ӿ����6�ˈ�ϻ���r&_�B�{��������|����X61�%����lv,U�f���ׯ'-̈́���x��y�+���hZ��X�E\:��d����P�q7�cǃZ��?S��.���w���r�GD���G����hey~�l�մ���so8g�)��+��/�`�����o����������]2�[&ưpy><)'�Po��	5��I�F��lm��-��?<���Z�7��E3f|�ЄRN���,�����w��.Lr=���/��~�&��{rK�GI�-���j�wj���J�����Z�!��n����p��g)%��8�ޓw�mY�tM���=p�kjz�e2#���	_��/boKm�3#���k���x[���N:w�|��=����a���P�~���~�3|��f��u|+tq{�a��[qX��_ 9�|l�����ױXo�g�yP��t�{��Cy���� f\ݸ��̉��ޫ�:�NߝJ���E2��B��q��;r�_���N�N���w����j�N�x�,4��:ߍS�g1���Vi���X;6�V/ϖ�iʐ�n���H)M� X+ZF��S�(O�*��Mf��w�Q����ebO�MX �Y�׬_�Å�H=��1;ϴGd�;�s����G�q��}�L<��q�n��_J�S��ĂM�al{���GI���8��xwD��2T�k@V�z�� Ώ�{���+���=�\���='�q�a�̳~����L5]t��n��#�6Gp�񿥍u��J��Jj˵<X |��Z@��'Z�z���\fPdn�L��\�a�� Uȕ:M���$4��I� �'��h|^��P]���Բm�������`$?�s�+���X�x0&�F�-T'��U��N�ͷ^�Rf�^�����.�0Tl�]*��oN�-��L�Ϫ�,I���R��%�Y�~��彯x;?3�����u�Z?P�$�Q5���3�(�'����0MV����h��-����[�Md��%��H���u����������P�^j���{��S��>R�
�z����%�Y��˻(.,���o��a]ו�����P]n�h���>�!�BY.��$v�~D�?f��V�3�ϱ'&<����v��C/P�,9�
�*[����zY����90"�C��˥���?���i1^���Mg�:����7��2_aU���g��(�j̖�|�������Og����kHR l�����J�9�o:��y2Q �|5'Q�kT;�mQ�7�IgJ%�hb�|!!�p`ĭ����*l��BuL��Ҧi���D �kA)<�k��x� ���j�`Z��+n�'h.Kϵ4ּ������D��P1��hB%.T[f���G��i��{�UՒL0��b!+�,�j��)�\  ����s���1�n�d�>烅@�9P6q.����Kp���P������I˳#���v����ͯ?���������6!���l�N�IF���H�_��E=_�u+d�㳲e�2P��=\0��[���mΞ���V\Cb��w�����<�\�wK�������2׃d��L�a'B<6��8�_0�Og_�2�,6�c��q��;>��c�. ��ٻ]k8$ ��x��U�>u�<UJ�ܭ���B?(wVq�I �����BX�{�vD`��fg.�2y�4ݪ��u60��>I�9��a�`.	Z����W����PΊF�f���w�z9?�$ىt+W�cE��Iv��?�����oߒ��4������A`����D�|�u�JUV�urJ����R�s�^e�x3��xt��������yi0�%�>Ƚa�K���z�H/W�o$M����v��������*�rY��Ɩ;:�Ҩ�*hW3��/��#�<��čЍ��j����������Bj1�U^	ƌM�޾B��=��T�5�#������l����B�Q�l;d�
sznq��A�q��=�F��E9Gܱ��`$͜e��yæs����o	�F'(כ�ŌvebqJ�.�M��~�ev��m�,���KD�Fu̴e�>�k��E�Bg:�ϸ7���RS+�sn�����u���L�СY�F������[�9����i�AG���e??_��2������a^��M:g��Pc�* ��Z�b��Ix��e]�؍���i��r�Gq�eCЯ�j��^��%�@	��=���;-{�[���u��\�H1�y¡�eŬ!��0l�`p!'g2�N�P�U���Hc��\!	r`�2@v��0��x�ɡ!��*9]���\��"�V\��7<�C�N�;�##�](H�Ĺr�â��KF$��KK\2@�(֌�Y��d#]qGC�L�������3!�,��F=��+j�N�Gi%λ7x�ǽ�������	ZA���T
��Z��ѹ� P ��_A����"j��IT��,iw���tc�l��?�1x+��W�Ǭ � ���pj��t��[t_.;�F̪ʣ�P��Q�h/����F���mOJ:Co����4��A�]�
���M�6��,K���rS#c<���@Ҍ��c���ı���O�/4G�E݁:;(/X�ٕֈl�Ia�����`��|��/^�/�_I�v-?�XM{�\����8[��|;�8{�b�@i�.wd�F����
��8t�ҧڗhR!���k�C��N�ߑ�7Ym�H�/0�[�6�eWׇq��j�uT��V�Z&ZN]lh�Rp�'�q�9d?W��41�?&`��JT��|Y���|>2�)�{0��Q�7�A��4�ؑ�ܭ�����-�V�%��H���bR.�F�?= ��/�^{����y�Y5!}�1����n��!z���w������+|x�u�ERf���
��On*����B�Z��L�!B6�G>�n��(�$�H�%\ ]�x�u	�2����)�]po�����sy\í�Pg7�[���� �R�0w�6���㣑����
�O$�d��$1c.�e�cx���.�1�zW��1U������(�`�3$X����X.�Z�w- ^E�J(+G���M������?M�rA��/m���띙O �Q���5"�Z��&p��Y��2�H8��)�_�� whI72����&�r�������e+�����nx���Y7Ȼ󕟑�׿�s��-)['�B1I���Ụ�6��D���)�ISw,R��*Tn$���8��{�������؏,֫�����u}�*�	�x����?rDϻ��ُ��D��o���"*� �A����Z�kֲ3�n9�Y�)�	��r�_?+��ڗ;T�K7/t�Eo���@����C�Ջ�4�˅'��?�9���5���Y`�Q��׻�Jfo����su�X$�L=��x�y��(�S�IM!AC ���,˕*�����F�vڊ�ó�n,���='�n���e�1An�z+���t��-��xG����%F���YD���Z'�0wZ?߉"�|�.Щ����Q���1xlL�/�ԋ�t��=6�[��τD5�C �K��!"C:i�D�$����5{&��aAz�@0�>�P�||<�w���~[iۯ6�#�7�s~}�����qJ�ŹR��o�ރ�����[���w��~�z=)����V�s�2�/��k"�e�A̾��|Oe�x�~b8�:Ã��O8:����D�p�j/%�3�y��ql�52�O��ے�n�D��u#������u`�(�V��9+�����8h/����8�-.=u�5��otK�
/�_
�h�^�px�+޶|��=6(�?^��#ى�*���7o>7 "��,s{���	)~�|�����!;��h&��F�����R-���l�rV���(���>ÎU덑` �:���^�Y2q�����BĹ�~πK�A�2ݳ��-�#Q�ʐ�~�M�n�5%��7�v?���;�����\�q���t��0��0x=��߆���ؒ��o�"8z�nWT�*����hC8C�W� �B��"��8���ϱ<�C[:�@�<{����A�'٣R#��%Т����k4�� �p��C��o���\g���}-�5�Q|=�O��z�@��5��)����&m�}f7rR�B!/h�������X�z=��b�i�:�>t�������i����17�X/���� Teд��Ig��}b���צ�$w�|]:�k���깈v���."�&aj�=	��F��h��O�b����w�7�?a)�1��<-BTx�����˹��͝`����,'?��1�v�u���+AF֯aٹ��N%�s���Gk�IQ�v"�4��Q��8�t!s���I��'�)Hcީ�Լ@KD��K���~S$k�Y��n��^@�_���vA�=�q�a�}�2����F��F5�N���bp�S\R�`���[��~��|�/�t( �}?ѿQn�V8�?! �O���L�~�Bx5�5�;MT>�VM�A'���{~�kީt��\�9�P;t����-Tx=�s�����|g��+l�|Gk?�Zo���i�P��T<��-N��q�=,m���'�A�ED8=4�߆��E��^����glv-������hjWw�`�h��(_L
Ps?4�zZ���S��v�!Ƙ���Ĭ�{�G���	��s�T���#9~�?n��i�z�o�%��z���%:�M�B ���-"=v�v>�W��<F�ӜZ(ڥ�Q���OE��2(9�J�Nʿ]q��>�B���#3���
!.$%n�T"��*�W N����g������|�[�]5��f�$G���;P[U��^	m뢱+ƌm{ƶ��m'3�mWlU�v*�mWl;���{�s�������xƛS|��M��ﾶ�a�X��2��|�L������?�@���ZE�@�9�|ܠ�_뢡�5U��|������HO�P�V��.�w�ʀ|B��ykZ�����0��N����~��j��lT���h0�GR�����%3�K�">8X� !T(vZ>su=o9u���;��Cn�Kϭ7N\Wv�v�~GK�v�X�L��'�;99kVf�����������,��p���W	����[]�.mVN��`����&2��5�_�G�d'҈����!�.J'@����p���'V����m���?$EI�u�7]��{������j2j��K��ع|�)9�8�BN?�u'�q�R��UL��ѽ�)W�C@)��?��:j��������S�ޔW�*��3�,$5��hD~v1z�H��dKQ�5�/��n���-z��Ci��H��(��)�����m��&}�	%U��M�F@eLB��ax��7�F��{���B�������`-N׬���{��?�}Ȍ��ѣ���ԁi5]��9��Q������<ִ)�h�V�o�W�U�}v�����([��T1ϓV�x�AC�faU,�Gs�|2"VI���5B ����nuBܡ8���y�����yz5rs�@��@R����sd��0ق-g2�i��?��Ji!�:�s�<'��4
�/B���'!:X$"0�����'�lԟ��.��kGP.�0�$������c�.9G����*$T֛vj��X�>�Θ"�%�6��|�+B�6���mY�	�߾���l��c����PD隿Ob���\�_�M��a����x@�F9���=eX��2Y͇������˪��Âa��O�n��~�3݅��>�^$RTdӥ����?�w׽�q�⟼��.0��t�ջ"�j��fշ�U�k`�x������&��R���
8~���`�,k��9�b�I�a��0-�h2��b���wǞ��v�#чw����/'b!��ϴ�xNw^��"��V#��͕��!���a��weTv��P
ӻc�e��QMY!�s*g��	M�Q'��$��4���S�q%l�js��x
��z�l�ό��Z�U�b�D6�j�WR��B�5o�ES�mvf�����Pߣ�d�$��-$��L�������M��Z%m��/<mC��$��T�+,��Z�"��9c�f��o����#�����7"^Qh3O��ґY妱Ẁ�f�.y"�>�v����: �>�P˾���Ʈs)�ܾ��N�^��ǖWD��F�4����֍:��ܺ:L�)+y�O�No���׮�G�&�����.Y�B-y6���w6���]\zNՠ�	)b?l,,,�M��������y\�T����_'V��j3�B�»u�5UR-�j�p~�F��F����Y<��z����E��s���e8���vMܫ.�)8��|ϧ5L��8f�{%��
�,��7N��ȱ���Yc;�*қ$4��)Lԫ0�%��A���T��Om�V
a�-�Q@Bv&-���KK�����Ј��*+�������pE�և�|�f�;K����O�#�Δ�\��������B�:u���RX�̬�G_���ot 9�u���b��<�N��i34j��OGgtDk)��:qu4c:��0+�*+n����ئA'�X���W�⾨G%h~N�K��)�ӱ���ۢF�#b�Thq����� v܀^[��}�4 y�@��B��K��+�+�*�
�I�5��KC|.rv�-7��Y~I���N�H pg!�ơިZ6[�i܈T�/nV���ۗ����ƻ�"�bU"�ٔ-��bC�Ѥz�L8�k 	1�V�\�Ϲ�������3����6��9��D�?�n7�&<�*k�Pkmv�E�u��PT��Q?ñɁ��`Y�b�CW
��U���𡢲�h�KMJf��Ji&��s�C6��C9DLSfЛ�C�ѹK�,2�B��Ol{�n���Z���bΆУ%��#���?y���.^��O���o���V�E�o���޺9��sىǯ��b[�ӏ���Fu#g�&��1�H���,(�$[�^B�������!��P�'W�܄.�Zi�b�R9�����㯢|<�&�ᜎ�̥���"�`�!�0��*�_'�I�泋�An!I�'s�-D��[��2��|p/�Ф�w�q��}��3�x*��x�a��Ҙ�x҆E������ثHٌH|6�Ы$���ƍ���#��c��+�WK������Ҍ�T_j{ƿ���i5�N;�w6�O˚�)�&�-iGmh<�C��@�:�<W�2������[�\�iyc2-�6�Qɕ[W¡? ��Nٶ�h��B�kL��]p�<��pm��m�"'�Tj����C�oW��4���1ql����F��C��**�\UѬ?r4V3s���'��Pk�C�R��Rg�]-\^�n�9�Ѭ�	5���^�%.������}��1�-�����8�2��}�
~������N�K�����O�"��P��Ow�j`����1G��%���j��u7y�
�	<|E+Q B�qձ�S�ġS_x������|�>o*{$�Z��x�՝X,Ofh�#���"�����`�d�XG�q뙊�v|M<�kgaW�*+1ut�;F@{ՠ�K����4��-�N5=wU/�.?�nˆ9��sK@��i���
��
�^�x�Ou�DR��5ّC,��a���+u�\0RP�DJJU�wm���&�L�ಅ	�\��b2���y���,A��k�~Rt��w��F����;g����_����	P��horh%UՕh�ز�5��t�V�	��q�l�K�)kT����O���sk�q(�CQF@��8>�~��Ȉ{�#p���S���lyL
�]�)�G��b�f8X^��@
��S΀߄XXH�J�a�u�5�����c��i�A���89|�
����F��`d4�R���bw)hX%��#�f�8�)R33��f��!I*A+�M"�;%��ċ<�!q��(~a6ElF��	ӈ�$�\�Φ=��޹���*[
����prf1`J��-���0�Pcqr�Sb&��Ip�;�1�χ�!IbG�Y~�P"���9���߭v���ۣ͟J��	�s������Uz�E����@�v�0e��)���2�o��N�8�[T��\Xb����A��^1*�~�v2j�
��!�O��Q�s����৭�dv��[xI^#�u�� R�d�y,<��G�=(�!��RRQ
+�eb6ƅ�����h�ޜ3�\aT��^��+�3�������|��Z�7~���_�ԃ�L�����Z�H�[� ~���\
9�M0�!2w1@�ì��[�
��gL֭Q���8�Z!��U�[���.��TULQ��9�4F��T,hr߹�nzW���Ã-��ԥ��Bi��IR�����ɜ8��;�<r�o.���߹���#�*w�ܜ�h;��� �JPL�B]}񟰰[k��ƈ�-�W�{��I�3�ʾ闫���;47ؓ${@�j3
�w6���+3�^%��U����^0�t{q���z�@�˓�b:���"�g�N�A�*W�Q�M�1*0�^�{8^@OV�R��>f)0�\�o�0dh��)�x������R$�w��y;Qc����\�yNɵ*��(*��'H#%Q^�7l�z�<'h��y��=K,�� �M[#=��ᔐ����<�d�҅��I  ���?��P~���~q�D$$��j��`��{< �Fn*������o�g
J���yޤ]�Z"A{���*��A�D]����W�/Si��!�������V{���HD�!�@pޖ҂^��; ���~�
�KC����+nT�ON*!">�ո���f��Y��$�$�HR�N��[S2Z�(�luᲰ^[�[��v]�,�&/-*Z�5}��]f*�u�U���(�Z)�4*��5�L�h1��Y���	q�w�+L$�k[٧�ޑ9��!i��䤔���@+��)��.&�O�v���FK�eGx0���8>\3�!�-3e�N5k��&��;��I�}t�k��<��B^9Z�Q��
I���i����DhH�o�ж�O�٩�&x�
i���s��~��è���6��"椠\1�Wm����;��F��#����eH�}�8��k���F�o<��2u'��s[[T�����A�k%)�_���d(靲M���+&��	}�J}q�1<��ú�s�oR�NR�&�f���˝�������KP�� �M��63��]��Y�%ϓ������4�A��LK���ʁ��0��w�<�o=�C�hK�ŕ��NC�x5%^�>a�_5z�(_p�=\�S܆1e���ϡuV_:��R��#ٕx�=��Z[w�P	59�x�0#W����uxP�Q��@ȱ�۞�x5m�t�߻?7]v88�9�5����tY\��*�c���BؕrC�kz$�P�<y~�6���dR��;���1���13¶�8�O�{�9��}8�� AULtή����v q]��8o�\��|p^)\u,����nzO(�<W&u�E�� �3�������H����2�**��B1f���:Y}�	b	� ޷#�'"���M�<�%c����U��I��؈E�`v�J`�d�Kʉ+�Z%��	�٭�Gd�(h�c"����W}���f>.�sn1}y��.֗�\qD�6��ק~V1�LXzo�y��0�TЗDho�uӅ��D>�>��7Y细'y���V�bˑ!J��K6��z���b�֯-}��>�@���;1T�Ç?	��/�uT�x2��a��5l=g��6�j���0��ݍFK�� �7��'U���T���Z�S��z�C Q0Q����a���^]�6���豜l_�Ӎ�l�08�Z�F���m�8[�Ȥ��^ѽ�H���o���f7��#ϸ��ݦj��/Q|;K�v<����%����py�8e�"k?��ܴ�Ϸq�C��*�/�����F%9[��ucO�������S�����.�u=���,Ĉ)��ڪ�$yj���%u�9�U�������Im�S���\�_��.��Y��3H9_k ��_�J�4�S�{�r����K�39���h�pO����W~�Efǆ�p��@��+��D�9C��BS���Df��~"�$\|���>l��c�J4e���yI	��h��~3���_,�Z&�� "����0#�Y�ʱ����\�ߴ]�'`�7ZDA'{[>�}Hq�N��ĵa$��WF�Pq����!z��vWZ1��f� ���߿�LO�2�_�]	+f�>}>�&IB� �X���ʡ�6�R�i^�׏�ްF����~���$���IӃU�Vuj��2�GM��F�q��4i{q�]��s$������M���Mb&�6�i��i��1~�,�S��yk�6=���Ţ)�IGh;K@��G{�!�|�=#�z�5�FߖT�U��,�:2��r��f����:�
@.�:���l�;N�e95�������<�w��h�Q�0T�ari+G>��54�Z��?|3��-RS�$h/���x��ܺl)�0�.i�8�ܠHB\	��'<�H}{������x�t��O��x�0��恣�P�1s R��/��d�ty"6��},5� ������{aw�/��T���������0�o�Or3WAOz2�D/Mn�)�E!uӪ����Pz��uAw5�:]"��n �/�'"�6 I�u���A��T"X�V�f��_���m1n�1�>xa�ԟ��r��Vچ䳉0A�[(�^!��?�̸�h"
R�:���(9�*./�����q��wJ&'�%ϟ�����&P�w�;��LQ�a<�U�-�=c�_���wp����U|'v%��=p�ƿޭ�./ni�0�kj�C�9����a�oJ�}L�ljm)��&��P�x2@�W��I����c3�%�)�*��5�)a#F���9�u��|�N�B[��ڱ�8�K���Uw�z�s��vM~W�TP��7�>�~�t�v"Zma`�B�{h�XR��� mlΖ,h՛q�{}�g � cY���m ��"��*"��E�S<FRBC������`�V�X�U��>���H��N�bWM7ז������-�b2�c+6������%"�{&�;e���|��b���$ſ��6����m�����{���X78�(���q��e'|20�f7Ny-���������U+��ࠉt;3�G�jMl��v��专��O�FO�h�����6�j�&a�t	=��k�.4~����].
{��+��Qm��4��X���.8b4?��|y���
3SD��J���q�R��(��5<�_i##��NZOb*_4�]�e/X4�#)�_Yi����n���ӐdZ��$Twn����=/��O�)��������3�e����ة:�{7�6c��e�$Br/�<�$�9�:m��_�"���}�����cY�Lt��y%��u<�{��DڗLC_�;h�k0�{P�ޟ�����ٳ>)������$�,�5*�Y������W�(Ǥ��?�
�U�H ����:C��M�8���\�\�$�ˊ��"��;����:?�HE?���&�zJ)��B���˫���춻�Y!$�J����ԕ���q/�N�o'�c�9�)� �x^E�(�:ur.�������!��ⅸ!C�j��d�l�Af�<�SI���HJ���#�J�^�X�3��ּ�1t~kpM�$�CVj��������d��Y|v��L6��D�j�;�Ɛr>���V��IO����5��3�����*�����)��o83_qN�e�������`������=���a�C*w���"��s�R�'���9��jx�Z�%N�'B�W4Y}Q� %�_�W���:ذ%� v�e�{��S?�P`۔���Fگ+� *B�&�g+Ds��m<�kd�b׀t��ӄ�c��5��rX��k���?���p�pg0�%.a�>7�����,Z[��� �J(,Y�R$k��R'aI�t��*���B;N�=�0Z��w^��1c_��d���ʻ׶��h*Ap��M��Nk�.�̖���;MX�k�ĸI�<�:K�vy��Qn�0۱� U��K?ׇV�#,`��	
R{���?Wku�DS�S�ґ��=��V��K$����,Z��(������K�:�ݮF�a�<?����0�C�e�Y����_�����A��=S��Xé�9�T)���B�\��?��M�=�&�K����9 ���T��Kg������e���Š{^�7��rD����)X�w��Ota��MH�nE�{"�"&C�r�����Z@��������F����E"���J�T �u��f�v�V�u�&��v�$�G� u��`g|�q=M"�G��t�ZΘ���}5��nau9E('&W��bF�\:��2t�̓Us������mA���5V���Х�@*9~�O�.Lk�9R4_���x�I2�^V�{���?*���4S� e`'	M��j�-�f�!ȱKU��y�!D�Y���j��.{	�"�$ޱ��/�"���"��1���~m�@��$�VA�\�W'��lG<���#7鿣�(�_G?eUyS&(��&����*�^ ��H��!����MJd����
D�B�5A�p'�#V���K�J�FR�P�
�T[�PA���\J��|?,����[��|�t���C��m�ѫ%��.��������'�Ĥ)��^���	2ˢC�Jօ��B꼑�[��uۀ����z��B���\ү!�9�+1���4�<P�\�su<�lNI,>�3߽ro��O�ayl��ۓE�����뿼�Ւ�� c�h�ѫ
U�rzLy�X)s�"/.!��Xׯ��8��t^y�=#~�&�t^w'�E$�{X�P�R&(eBn ��6�D+)(�����2[��O�M�pi�RX^�9"��87|t�N�Ц�x�#���׶߷_�!�8ԓ�N��"�M�y��0��-�_YY��8e!e��I�Rnnn1�{ʧ�u��AA�����h�H^G9�,>�=��Q1P��*�+9��/���&|�Z�2��zq=�/��KhN���2��
�	�����TQOx��Tl�Ca��Q�R��q�eF(��o��/O �T=ڗJ<�O����F}v`�L�E��WMm���X�t+ϓfo~vH�9}��륊ɹ������O~��iɱ����x�W�5?�M��L��>�nTo���1��pu��ƄuƦ3f%V��xsE�Q<<q��a��su�����s1��)�6��.3�
2'�gup��wq��>�����IufC�v��g��g���V�{���`[+��zeAkG"�b��EI-���i`�t�o�a	������P��˅R��V�ur����R1n�yQMFP�t{�@����w9�o���>'�����}XQ�{I]�����g�o�|�b:���Gt}�p�C��{�l�Q�w'�1�m���n�>J�Ԥ�i�{y<�2��UQ�� �Vfz��f��@���ڏ���Q�)����5� ��90
���w�#�#����n������RQdB�I �n3�Lϓ x����7��e���"����M޷Ӥ�F�
���A���s	�]������x4�8r��3�v��0�����2�-��|� ��FEJ�}��^�����^Y��H�O��~Zx�jKi�<7�S\U����sg��};.W�fĪ�	ކ&m8�����Ҫ�S��U3M��Kě`�b�k�_݇�N.��r#QǷ�v?m�b�/�i= �F�]{��8��;(q��#]ʑ"�u���8c+��րFЂ���:tLAY���o�Qd���_����ڹ?c9�n���Dq~*�M2�aZ3̏��, 3g���J��ޘ�c�>�QٳCq4]�"���:�Ǉ��"l�k���=�^R���<a��<�2&���$���!�]��>[+Au(\�#�۷�\c0׃I�fo�M��
Q�&S�A�xZ�D�����,�@�]X f��G�֪x�V%���m~����
��t�;�ðH����pӁ�,��������U��uD�njMW�O��7�]�ru_����(��?ö�9��	��>�����f�<ѤN7x�r�Q!e��X/Ut��nK�]�ə1F�dF7 vi��1ei��wU�Dy@+�j��e�{���&Lcs�p�qa���ͬ�j�=~2��_�f��f1��gdJ����۝�]�����nw)�l�N+"b��f�[��h�@�`��wN��Ch��� �C������a!���b{!�J6��03d�:6�憎͔���b���'K������Q�z�uD�?Q�Z�A���T������>m�����ovm.\� Wf���q�_�~/.@ILLL(�'������/�?� ��z�ee���#^��3B������5�eN�ک�����sp�NdY5�$Wp���w����Ocr��ЭtI�V�\2xU߹~v��ф���҂F8{�kY7\9�qu��:]4	3�H���2i9�}~�	V�3-�*�'(�_I���h��������ذ=(p����//�ЛZYGo�s�ż����f�Α�(X@LXcS�P�6�JTeN���Sﶾp���ąp�_%�VI2b���o0��9qZ:��5�Cu����Q��~b�M*�i�&�3Y�|X�Aƌ��G�����`�سu}|�]?w�_�,�;V��ȁ�7�y|ꔦ���Ѡ̔r9��b��-��Ӏ��*��	 �<C/|ss�M2hR�,�,��T�K�׉K]}ѯT�l�9\�ؓߒ@,��#^|���޸�x�օ؜��cC��_��Z�/v?n��w¸�{댋g��UjT�@���/�w����`aV�6��Xq�P�hO�O~<��򚂋~�\z���z��B� �5����(��Dc��P�N�V�p��[�����T��u��%���{��9�s������L c�����p��f�ږ���Ě�&��D���b�D0���`T��0Q�oa�.���moS9T�-.��Р8M�4�<�ƛ�s7O&k��S
��&��e���~sFC>*E�F=�����I�Ō�-�b�W�2Ӄ����RA�|��]����q����q9���4M��T5Q��w͇�Df�'uI��1h/��(C���q�e���8-�[~�ٶ �0�OAW��	I��`4&;w��fL���n�AY���O�~]���7���n��MZ�[d]�"�����\k�Cӫ��hJ�4 [w3gR�3�:3gk4^5�q</fX��)���/�p�t��
:��j.hA|�z~sA
U�R�_�N�1�?:��O��)QSKW<��E����ٽ��s�bW��k�#_DJ��~j���$i�c�֚=�3�@��xa$�zw��	����:(X�:b��!��=�ݒn�bjٜ�'��˼�o���6g��`��	����ـCҩ���F�ƣX/�֣&����pb �I����@d���T7iVb5@;���=�P��?�ע\���ce,Q1��l鋜
�Tм�h3�rݢ��ߖ�e��������P}Ӛ�B��%�E��ӹ#�P�ޮ����ј\�$��x���;�7Ў� �sɳ�`aZ�ؘ����{eA�s�STY�|��CxcY�0���{�F����j����^��Tm2s-���>߼��R�^��ZxT����̆"�|�L�5eg$\$Я�/'`���\,�Á|��%Sr�\�9�c��L>��M�F�y6�ՠ���R�?�c�WFط�����7��Cb���zrI�L��$4�"~�Ӿq�!;�b�`�Pl�I�
?����3:�EYJ�b�U��v�PaI���%���r�.o:��0�ʥ�=W���y���v�F��*ٵ������Xo��a��p�Z��p�@%\��]��$^�����\~1�-fB8"980w(�*Ͻ�����+2�i�ީ]�y�<<HY9�<QQb�6��_&+AD<lÑj�.:��6Wra�tL����F[2��e�������fikf\%�ݱ�MM�,!/�<wEj�݉�k*e����R�1~4t�q���r�~dfh��mr���=��o���Y�^0_A�RWz	S�cI'niYtﱅW��������A�8� �c����!�j�W&���e��(b^�Ӝ�l�{�zx�ղ�r,�OPav��*�}B�r
��U�C+b�S�q/?��k4�_y����h?`	�L��wW|~|D���ώ�c�tﮝ{��{��B+�߬�zG����f� �DFQ��j�G`d6�Y2Q�FD)��9TĦ6N�� ����f����_�|6v��;��=�A� ݡ�[�f[��QTX�"���RaY�~���D���H8�'Ӱ��NCS@&�o��ľ�/�i��G�5Y�)��O��7g��l?	�f4���~nr��K��0^�Q�d��e��^ 	C���.KP�m�F)��� ˂�0Cf��,����C�V�M�T���;�b�^:У��A\��X;�Q�6� ]��pÆ���Q�נ��lʎ��P��y	*����u4z(�Ŋ��5�+dR=[Af�ɑ1fp�}���r~_z{�d�z��ԃ��*4ٺ�	�>�O�Ʌ����4�K~�݅||b�j��g��C�O#����Н��Ϲ�"T�Q���J߼�^�|��5Bd3Um�"��T�=y6� ����S��	[�^T�k�Cˈ4���m4����SY�������n��t<]��3*�v(�J��À:�5���C�+��9�Jfan�20�37�=e���`͠�K~�%�z�֦Y{�K��^��~��j�ϪNzĈ.������B[���"q�2Dfz�����d�����4%����*�ɡ�2�AyIw�i�Ą0��vy�"l*�#�CuE�Ei:�\0�+�9�K���E�]������ܰ��q4��!ҁ��'���K������u�:P����$(����XB���T@�$C��XP�pn�߽��ȃ	�����h�ᯋ��E,º�o�ָ�#V��c��I�? �?W_��y�f���h6���?E�2t����@��3��z~dB���$+{���X9�aE�#�؅�W�wo!�k����tݐj$�%���0ęo�7jLhn�@�����W�fN�C"y�ot+���b�_��T��|�L�(�S
�@F�a廩cBRti��3��rp��@nU=�Q��˼���DЬ+Iv���n%�3�ʫ\��R� *`d�dzة,G6��V#k��jA+�&*�����e>��C*ܤӳb�,��n������h�ՠ(�h�Ď��x2��2���1h~~������4aw���G�~����3*"ʯ4/�Y�(p�v�� *�{w�B���+^����^��ո0Dx���7Y��?TJR1鑍	9^{�EָǶ�Ǣhؓb���hj5��?���4:*��**9d������^�f���3��8s1�I��x�>-B��ʿ���_8mfC&VUJ㾙ε�;��a�/���g�TΉ)�q@_4���"����G-LpK��؇@@
\� M��L��C���#�:�-�ɬWR�/�V�Y$t�n����#|��d|G�@!��2�ޤ�XCt�HpdO%���;9��h���h�4b�e�0р�NU�9sL�f��6��e�Ӻ��\w��tgp�K��z��-h$7aoA{ ���]�d�L�
�#Zʈ'��ORE��tso�͸��m٘���B`��S�Q�՜�/��rE�v���������j�])2���q{:}y]+��l}!� ���5�l����Ν���X,���^�0�)g�$%�50��҄�iͤ(b�?�)b�/�IHW�ʷٕ���9�~Hֻ?�Lw��q�����<��V�(����;�����w�=2\:�2i��+�F_|��M��þh�PH�3��7'3�F��)�+1��ŨU��O���½� |W��O��X��if��sMh�G��액^�J>j ����<O�I�_Ip�IZ����w8���%��l�$m���AW��\����%��8O����//�/#������z?�eN�c{��S�����QL>�Yyzm�v���e}��j�Vӹ}J�7V�G�e���,/�4o�E�dD�F�K<.7��d~�H�D��ұQ#*�YY��NM������V��z(�KQ�1%�C/���N��S9h��{��YL��R�aP���*�Y- ���P[V;�`$�|�8��""�4R��)h���/bY��ݨ��hi��Gܫ�v��F�M^�fx��~.M��wK.�x�험����[NF�	�d2�i!�:�[!��Y�,���\��u�Ν.F���_�ۢ�8�㻝��`}o��}Cl�
�;/���s$O_R-��He#��	�a8:��y˓h��9�HL��ūr�������<>��X�^����� �ݝ���ޡ~Q��	�� ����˶���5�x�W�H4�6�f��>�a����H�K^��v��>5�B�M,�|�Rf��ɺ��Z7^�6�:�h�5`�bO��s��U��y�iYj��v�L���I(�{ǃ��\Ö1-G��{�p(,V� �A\�C�^�ͧb���i�\�G{4z$a?��Q V���2�Ys~$!T%�/������s?��iغ<&À"痳�zHD�6'gZ�9���a��.��L;����;�po ᯤԆA��/�~5돷������ŀ�g�^��Kg��	���;B� �(�o3v9�dO�S1ͺ�F�K"�ly|a�^1�nR�}Jv��uB �Xj޷��FT�����K�4� �$��	�N���/i��������H 4^�vD�c�R��u�V�=ʔ����H����ו��X)���(S��)[������
��du]���㊶�"�q{���� ��+�3G��v��Cy��>�[��y^��zj�񈭈�\�GG;j��K��7�'�;W��a50B����k6A����>V&�׎��.�$�/��>j2��M�����J�ݞ��鶹l�@�4i�p�t�Kc���r�Z�/��h��cmÆ�������2ӱ-���F��L�
;^*a�*'�a����޴}��1rxv����y ]:+$ig��Z����O�u9��O�,��?�T�cH�o���(Ǉ��$S���p�0NǗ�>�IAc�)����䲥	
)����;��3���Xx(?�ˎa���'{0+F�a�b�FMl�R[�%�Es��q?ݻ�@�0�	����}�}	t��m��"��P�ˏ$.��;i�$�Z��)�l�b4�7�^Va�B/w��v�Y�w��jԌ��(F�S "��B�P��R9^�a��+��Y��|�M�5���,��eR�ݖ� �\��&o��Q����#��9!wl:}�i��^t��#׳���ͽ�+�Q���(�|���	7:Q$J0=n�p
�����d4�=�O��o���.KAk��ξ��l�S��æ��&PoO���r�usZ(��8��M��^=���A� zܶ�Q�zNC��L����Dh$,�q,6Dh�QQ%Ҳ#�F���D������툪UÏg��߆P�?�%(+{-�!�b�LP���Y���$�>��Jf�bʕ���Fr��&2ב��i�0�b8�+!��k�RF	IR��C6|��"A�]�5����
�3���)C$������
�;��i�]�͇�.$Zy��u��_]e�3lƂ�	#�3���v�Y�bxN=�n5I��4�ĺ��s�+N��m�E���#���g�B���I��?mگ���5M�ī�,���]%1:���0h��`��9ܪ�e��>�����Xf;��9�"��4�ӋZ�/;��}���X�V�\����ONlF�[�����s{�P�}�=��+k����f�V�=�4�c��p����6@'{!�K�c��3������2nry�!#�~ݫ� �;�&�G��{����Z��3�L�%���r��ÙM�V�.|��h�2tP�֦�1/xv.㏩�5�)b��2��3e�Ҷ.���1fo�"㏖�2��T���V1��m����d�q\;��&V�����~Ӏ��+�����Ϳ�地�=>�/E�g)�U �-ЪMs	�E�'o��̎ �^����5*Q32�e�M���a�<B"u���k��f�M?=�q���Ǹ�\��ѱ���hEN����Y�\�6(����N��*�1L5E#t���ЍR&%B��	��7d�T�8Y�rpN�,��Ѻ�]d�e�ֈ�Ө��s����|��z_L��v��v����nT��o��%S�L�����*���t:H�M	��4@����|�s]#��ۜ�4]:sWv�K�m�Z����
V����BJ���@^%<�w��}x������a��y_�U�n��ֻ�9�n�C�|ܭ�q�RRXf�MҴ�q���d����?0�EK�E=��M��q9|�)6��^=�"��Z��Wj:��h��ה�ZN�K ��Cԣ��D�����>�:o�cf��G����7�[L���|�����W۱�r�M�PD���?m�:x�W�P�p�����OC#}�B��)e�y�IB����Nl;5������'��&(+r ,~׋�Mc�/?B H�jB���A�Z�m��}n%�GG�
�����
n$s�j���E�e׫H7Y"(�ŀRxi�j���X����]v��<�1Co���~r��))\~�t�@�Q��~�$ 3��E�p 5:₞�r,n[�	K�G�ʖ��V����$!Dm�z�K�$�z�c���Zsı��%�+�d\��.���ui�U�.�NDٰ����j˩��Ø�x�
�p������H�e�Mh:�[�d�l�:bݗ��,�v���zҿ��3�+���p��J�u7��01��(v�}�����A��|�U���e���	�yr�c2z��yP-}+�4"(������������u�w��M~{q�q���I�~1X��W��A��z��Ѝ�x\#��w���c��*���:��dۓm��d�6'۶'��m��&۶��~�����~{�Z{_�ot���������Za���;����3�ӫ�i�v�����Lg7��4�3ݹ���H�[�	�u�$�'��J��YK:p��&�����!y;��?������`�8�>R��� Dv��L�<��'���U�Og�-�c��߮?��'Qt[",��&d����b��Ɵ�T��}��5��Z qK��J������Br���)]�DKNkߘ�{�g�L��e���V8hӘh�����*����a�������N$��1w�Z�M�.އ3�+^�)��>0�Fe�+�[��uj lm瑩�V��ׯզ6��tNخ���c%��2{�	
U��OS<��.`z��Vdp����*Q��9��a��l��Ť�1�}�@�*�s�w;����~8��-V0|3�Q���,}�M�91�x�������e�^(�J���uTs<� ���{+��&~�� �r����P�<��U���f
�z�>��h���a�z*�Zͭ�i��L��i����j;���Mshf����k���Q�"$\�v�)�o��HN~]�~+�D4�?l�����b����H<����K�i�A�b=U�s�B�Q� �+��(��:�FIDq��YS��~�9�# _��q���Q	�����õ�>��=�=n���C�)�w~RU�&�/cs3�ؿn��#�:O`l�,fƂ���2k��_� z��w��M��u����^�pD<�u��eΗ�P&�3�\n�N���vY��}�9���a3��dcB�pޔ�N�����%M����3RJ��0���<.Fi�B��jQ�S�S%���b�w������'" ,�&�P��Kɔ���j_���DF+��ʁ3��G�0�Kh�)�٦ؓ�/��6	�����ǀ�Ǫ3��|�[hk�1���V.P��R���E�$Sx��	(�{��˘�푇-������ a@:l�i�W�^e�������N�"|��O�� �ﰇe�v���?����ͫ��IGiR?�'��Ɠ�nt������2�W�R5�g� ��S4o�I�������n\�ňR`[,X��6�GC�''1��Q��e8�}��X�8��{�92N6;�`�a(�y����6��F��ˆ�&M�nxJ`���\�_o���;KK�]��*���Z�d���M�p=_Q `�_�!���+�tͥ�ǸE(�8X�$%�$�G?��z����*�8�a]�G͏GN����
܀��WԵWT��A�s�f��l�Rj�����c���*#f�����"�_)�Y���C�0qjR��qh�m�Zm8���� �p/%�'�����U#.ߞ���_olxRo �̡����!Q$f�2m� M��+*Q*�e#�V�(��S�o���3R(\1!����4Vr�DΨ�-���6ςO��>�[����aG�2��&��`k�b7!�瓖�,od�q�hw���NԤ��
k���7��J)�U´9�r�)�r"yj�J9ݻS�r���� �,��q�����[f%�&���Xo�����6�!-�7C���cqIh�<o��_��Ѯ�=�f�U)K�L����l�'��U8�䤩��ٿ�s �����7��f������V�4�$�&�V����<�Ak2B�$�� �p����wn���k9 ���6��w�U %6�K�V�?��Iz�l:W�`��-���,O�,e6x�e�v��7��I��t;�_���,�`/I6~X-]/���չ��K�ӧX5y7�|�R �D]۠���Q24/�a�d���o�R����DΨ�h�L��nܫV<�˲0��W�񣦼�5w0�V������,	�2��z���f��n|���"R��<G�ަ�%ü"|(!ÕX��O�{��� �.��?�O5y�rs�B��Aqj������Wư#@ݛ��[2�3h��� ET�laO4u<�&�9��s���v�W�������g�B��Ц�nnn,X�p;+�z���K�_e�,d}�\,k"�4��ׄ?��ٔ,�C��V��T:���w88��ңM�)��OZO�Qߗ-�<nY��Pw]Vcs�$ˈA4���V�2��_K�=��B��]Â�޾�)��pr:�B��0����'��}=j׺�n�p�7l0�**Y��_ݚRbj�NTѓ�j'|]�MU�E�خ����s����x���ёM� ������TEM4����}M��*6mcVY㡓�_��X�^2�d�Y�HX��O��?�0p4I1�?J���H�S�0%gO�ձC�\~ױK�"���(:&j#�5��V�6J�>��/�^�&�u��s��7,g��/Y��,��|.��'*D,(]��`�
M`��%?e=M�z˦3w�O�E���[���|D�j$%<�?��ى��JELN1eE�4����"a>2%W?����_�bZ������nK��Hv���LĮ9�t�c�8��F�:mV���Fp2i\>����C���1a�S����#{P�?���g�VDv����!q�<`NL���t�xi��*���Õ�hTe�c�KDu�,]9y  -��3��렠�Z���l�ŕ*���Vk���^gI����.��Q�&��[�h��k�=��( aύ����y�!�M5|��ʟ��I��C��T�yw�s=�I�Ci6�Z��%��֯qo�p/(���ܯ��� f���[ßa���ĭ�;y?��+��+�$0k=ã�.�yriio5Ht�M@���<�����i�&��Nd�7{gY�!/��� ��UY:�zs=����=��]���_T2�Sd�d7,���-�N�-c���xzn�C��!��q������SB6T��>}��F�fR��AkD�T������
 ����PX�lǵ*
F*.T�!A���d9�:W�6�\��Q�~X�<�l������o��,f�����#��3���`cؤEF�NI<�����@h�ʛ60C��.�
.�)
[��j����	ש@�����_	�e��+�E�Y~��v�+�hZ���?��E�A����#aݲ�+�<��Ǒ�&���uX�y�UR��uD�Pi��9G��}�e����%S�AY���گ�Y¡r��̧��~�訶Ps�TuY_CpN���j��[���&� ���$"���wc�<Po�eB~ ���d��[w��)f��r+���J D@S����4Ӈ՟�O�0�J��K��gCvl�@�{��w��������HV#�e�t�7��'<����!5؄����/��P��s�d
�
.��U���va-_pQ<�j �E��c����/�O��>���=�!����o{9<�t�FZ|Jw^��g�N�ʹ#�2�B]E�Ǹ8�p���7( c�is~H�e�N���q�;��ۋ.�Rl�_�a���3�רGxe�L��ԖW�vCU�7���t����"���q+�]�֍��i��m�FS3�a+�������r����M��՞�-I�������v����Ps�a��E[<��0�+^���"�e'8��j�@�p�� ��ѭ��oaQ��/9ZG� v٘�&�1��R�K�����	�Ǎ�p<d�᛽h�����r�/�D W�VD�S���î��?����ê�:2�$T��Q�wZ�n�����j�D�$ѱ�pO�<��Ô�nI�pA��|�bA���計�P�y-e&W� *��Я���1m���ɷ���<��o��-�|KX�(��uAQ��5�`��A��bv��9�VX�ep�$4 Wo�����/l��y͂��S������Mϒ֊�P��m
#�1���DKS�����^E�Q׵�
�-��s|3V#���%��&��WT��66�[DD�O<zC�r�5"GȌ�wo!2nr^�\�V��@�w�~�P�����'"`̎9�,��1e��Å�ӺM/����?	�0�����D ~�V\E���n�YK�7���p�l.!z��tY	�a� � {o{
�к�N9��*��! ���v��݀�5������{����d5�����r��� ����i�i����c/�����񮰴��S+鐾�K6�禱7����=U�U��c�@�|�э<�8�:<���p��8Օ�����3�����U�c���{ �����L�=���ٷ��/'H�W"�4�"��ȯ>�����uOCC7lQ�s�a#��"v(�i�Ǉ�2���~7!&~>GRO��������R�m � ^p3q���h?ֿ[����v�[�o�����+�wij���<Ʋ>?�g�`/W,�56��y�TKџ?Z�Ѵ���.b?c��zS����u�0�V4�\��U!�ѡ�֐�V���6`�[�l�pD�T��b��<!�xk���k�o'�?�׏_k�%Y�j� z���7q5f���7jЦu������i�(���S
�������?� aw����:�\f��NGh���mHh�`�f�PG��_i�1q�O��g�9=�C��A�j m��)7~ѭ�sC���\S�*�e�P�8��|��5x�:
�\F�$n"���׍��K�|Mo&��c&��s�D�.M�#��֛�G8v'A0��3-�4�JK�쏥��%]�G��ۄ,
�,�'�o���"�_�'Ho��h��${
���!�G0���|���p���6���R8�*]_����,��j,��'�Dv �"vL�fB6��t�� �_�8�+_X���W=p�k�\r��W���o< J�����z�K���O�ޡ/Sr>���׾覄#����N�����N��N��*���쩇c,���mj��{(�cE�&�;�DZya�r�@�d���TK��@iʜXVE��{�h��F�E�l�����典N�iܮ��h��K1�����y_�-�ox<�@��y�Ļ$��&nl�fmEr2�A�C)U��T�$�h��������@���|Z "�u�H�u����6C�[�{�<՛-�帅��G�}_A(���&1��,�����?��.ᰱ��%r��h�wsss�n�tYZ-�z�|��sv�=�q V���Cf%2��<�� e��ö�OΊ���LS��Y�#��W厙���n���}�LI��6��0X�W�2�%�n{vu��������,�5����Xz�^�ynr�&N,��t'�x�e<�h�Z�z�����JXp��i�PR�:�!x���Jk���=�7'=�:L+(j!��w�����?u��ڪs�!�\Cr\��t����+��% G�7�z�.�e@��J���)n�.���a��f��M#ܣ��µ�vm�D����z_���A�u��|$ �vC�㻟㲋�G��fv�!�@��(��Ŀ"�� 4~�BZX��#��4� 	!�b�DV&��>�\�ϫnE�^~��w���{/�в���-�Y��~�C��bf�(F�o���6�-줆��+P�s^�O%��w(\�����H�#��k��Z��Ɵ�Ē�Lb��/�5��xC9�Ms��_�5)���2"�-/s⚝-�tƅ�M��^���̡x���3KW�}����wԣ�˩�N��t	ϴ�}7�0��s���C1��w ���B��=I���!�n��NT���א'ćE�"[[��Ԅ�!u�K�H�P���uJ��|rb�'�w�u������0��6Pg����<f~y]���o�e9p�R����|z^�7�'�W[�C5�C[�3��UC}����,8Ďg�8��OOk;��3���R�N�tж�RWNw=z�����f��$ٴ3qG?M����9-~b�xY��� ���&K!鎛L���nNz��;w�MlԂ�]s��X'R�l yr�*��¯E���-Ҟ�al.�������K��߁�l�P���&��u�8~�O*};�
5�/�tƥ������h��	r�P���g�e�� %�wF��W
V36�`0Y"��B<a �i5��c�;�)Þ����2��灥xG�;"���KyJv��7y��
��z�m!��ɣ6����#:ڭy��v�H�A0)�E�Ϗ���W��Ðr&�눛�׭.���?�(/��M:o�g}��T�t#�Xc�Z3�4�Bm�=
�eJ�ٙ%
�¬�%GK��K��T��Ի#?�C����b�{s�N4nw�Ie]\�/{�@�0��0r�ž鲐��+���
t���E�Q( #x �K��r���8~L�O�o"ٜ��]�cX�A��4ڷ~�C:�N�} �׶t�[+i&�N�l�H�׮�v�=�zw�%頩a�~������]���-�uۯ�K1A�EV.� ]�g$�������{|��^�jU�H�67��<˰�ȅa�V�x�~���q?�˔E|��.]@���������x�z�yȕŔ��I����}-�z�iH
(#2 �����C�<�وa4׻)TT�F�M��7�U�]�m���d;���4���5���{���D��žE�w0 ����*b6�L�ۋ��ǘ]�k�ԱO��q�I��~�N���»aoY��=N}���=�l��ge�Q/�Aۗ���0�ނ,� }�L�W�g��x�dY,c����$�*����eMRQ.~�nk�T�!xС�����?�f�eo�e�����㢗phQ�Wj�n��>���a��w��%���0�zhI|��JpZ.�5�4�%(<�D��{$�q?�1x��Tb�|��Tԍ+��b�{�"2t���x�:�9ΒR���Ԡs	W��UJ�y<^x{��ߎ�$X�ב � gT�h�AZ�v7:@�.k��f�T�Ж��-0���+ R������U�`ԫBϑ������yd���K.�*�dt���v��͙wW���svb�I���\k6�/��Zu�����n���1�!�#o|�`xk�m���O�@ $��_P������8^�Η��fB?9�Q��F���/���ս%"�R��Դ{�GG�{ʱcD7�v@�H,%�\|3�$#4��)���-�������I `�I	������>G>o����i�o(�܅0ӧZJ<�]�c�#e�#@g����T�m
]�!0�M�Y���s�t�搹�β�$�����S������g.K;,�	�'����)5���ۦ��m^��N��͌Gn��"�|W��g�WU(�׋?�c��� $���ȭ�Q�h��4�8 ʠ�T�����C>����E��#�pD�	���J����r�*�c�9A����7Y��d�i��͟��h\�� ��{��Rg��s�
�t�I�:��lUfl�_���<�O�2�����˪!�
�3p�K v,�j�d�R������zA`{Ra�Fߓ^�ʿ��.
Jg�8p�d��~� @���G�M�#�s(����1�����^[�/{dD"tl��j�ۧ�#_�Q,1�M��aĚ�<X�t|G�{g�����S��k�Z�t���笮�6`°9�O���J�MX9f�K���\� �Ƭ������(�ɲv�z#��BF5�����"G��[��~�=���b�v�~r��8d(3�W����y;�ryem��� >*��F5�E��U�k�Һ�W2+�MR����>��P��V��qJ���M��=��Xm�G�H@}y��4 ���|*��Yi��,��д��g����o��$���ü�#j�����	M��=.B��������qs�������5��v��O�'���U��#m�V���3zh�G����t�1�i�&�w���6c�Z��uoPq>���O�b&�|�Sp���F/r/���$��:�Ў.�f�%xi�_A�y��9^4+v.��u]O�N�%��>�ç�^H��?W�4�͡k���<8|qٺ�C�n&u���U� U4� ܇���C���������"ͯ��ϧ����F���sY~~����Ɍ�B@�lzGĥ���Y�ط?�0��9��^�8�)�9L#�����ly�`.�{Ǉah����b�x_�y�<�d�S�;�
7���~�����aᇐ����8����E��/��䰋y��q% j&�|��*�VyS�.Q����syU��dDA/S�P`i��ʨ��[�Br����`��餲�
�+
����P�P_����pT�,䦄W%T�DARQ"P�[�,`j�J��05Դl�!���(��E`�w����+��6��i�������M�VwM��J�X��\S8�\�a����ZK_��1Wd��zl�\�Vmiғ�$#��/n�/
V]v��Ȁ~~&v���̿b�f��u�Z�����1��a�Ŵ7N���}���3��9 ������`��4,	U����̲u�\��w������	9�	i/�e�yC��H���DQTэ�D�a�c���oWR=�^yv!���a^��LE��3�g͢sy=v+�F�\�>i9w$���b������[쳇04�qb]�Wo��b}_������?��(���^��7�����$�4�����*T�N�x�.�cܙ����Eg5�^{ؕ|���h������k��$��H�!l1��
ik�8�@ThX�f9�\o�&9978Oˑ�+��~���=�Z����>�&hp����j|�i�;13�� �Z/�7��{%�6di_�%$�<����o�(��u�S�Y�Ҥ�!A�i��SF��_��l��.��4˔A����zr8�dj5i�:n[��#W�+h-���#���,"����&ڢ���|��jt!Rմ��3����H������*��9��;t=
9W%7�1��hy�r;�r�E�**��u�3�R��v}7����f�5����n
�gw�6�vk�/m�W��"��摓6�����n�j��Gy�;��$�M������(1~�&�!���S��A�{0��9���*ą�	�{/���H [�M��ԽC�Tj�3�Q����4�r�9O�n�
.�qQ������Ex"�����B_�Dd�ԨY�II���Yf��d�E��c"�֣%�vF�~���	,!��o��4a�h�S��9�������o���S�7f���*���.� ��H�z?��S;ȅy[Dѻ�|�q��w��?��d$)�@��y��9����?D�Jd<�1|g'�e�	l�\�,��G$��紟'��zd����DC��BGx�_��u@��B
�2��Y%�.ȡ���j�]F^�T�/�O
|i= <���)�R��';��QJ@����-�ڂ
U���f�^�n�?�Hz$����Y��J�A���Z��W$%�gM�x�?��
���=綹ц���)�u�M��J��R��~��`�"�C�p
���������*�GGk��.K�i���"M+�cQ<4&�hxL���R��_��Ye�/��כ]�n��ӄ��SA0�m��/�b�ʭHC�Aq�f8���1,o�`Ī�aj�px��0ݰ��.�;o�0�P���.��pM���Բ��υYB�Ms����Ѹ� O��g�E�Ɲ�Ck�L�a���i��*w��w�^��s �Z$�1��'��~q��lPN���U�ƣoA���������:R��J�vАQ9)-g��b*#@�W����8#?p�g�f<>��/H��b�5Ǵ�z��f7+���
�й�6i\��v��?#ߌ�>N2? L�	MC�\b@���fa#0�h'@Vk�Wq�51�R]m|�����rYBu�F����4� �!4ǘ'�/֡�p��w����[p2�lɀSoIX���Z���PW���PΓ{�SM�JP�hѮa��N��r'�?�]^p��̄M��"��������=̼����5a\����� /oOS$v"sD�p��B7�v��x�a�����>�ćG��)M�7�3���r����N6��Tw�t�:p��g�}�u�.��"��p4B����
�
�$h�S��ryn}�4�����-p2���ً�zy����QJ7�ؐ��Oz<���&<z ��9�h�\�(����?�>�9͖��#'��$N����ʇ�glg�4�w�0����&ݴ���I!2�`��J�)&j�vqC�����MX���+�N�VG���b̫Ԛ]Y�3q�J�i��Y8�Tk�d��:�66��P�1����E1��q0�!'�d������"Ҫ���;�+�����A�Q�x����������	_�(O��`/�G2���[���!$KLU�9c�e����v,p-��|ɂ���nM��0��fH�Է�T �J���C#p�`����t�i.]�hh������<��HZ�,�G
A`��-@H���%(�����.V�Ɉ�;5��"Nk�*;��i����%��Iȁ��� �{ͩ4 ݔ���y���� ��|گ���|p9�|�d�� "����X
�bT/k��T�,Rdf��L��v���2���(�#�� �U�;��L��<���W&?pgbAF��^1:�ӨC�GH����{1L��63���Tٟ���x7�C�5�#����N�r%�-vh@�y��Ɲ���$��Zˢ˺��4�9����7gڐ���T�rhm�����+�.���2+ �i�p��
���Yj����i��ܦH6<�����K���Ŏ���2�-����Mؚ��k�J��92�g-�PI�����������%�9�R�A����}�`�7��WV�T��*V�͆YI��L'}�� �S�ԫD������F��L�A��Y]�\r(�# 	>�e�����С�c��U��rU��^�=,OЬ������lV$��kv'g�L�z�-�x	D��~3�}���p(+�nȁW��N�U[��Ӳ(l���%���k�}nA(|\U��KK��"�@���N�;��Տv��ً��?�ZN>��-�$�p�1Ta4!����7X9��_h�Cf/���!���{��-�NR}ևW�n�e�B~�O�Y��ľY��=��H��0JV(	��(�SÕjU�Wkǻ��_8�"0��Q��q[�lw��%Pq<G�j��80����[8�͒�VяM�?,�\z��hBoЖva8���n;�����G��:;�u��*����2?��G�B�ʘc#g�xN�q���d��g|lL$q���y?�BC	�H�����3w�>
r�t6��45��6��w�����2�^hU�ml��Ȝ1�����̆�R�a�+��\� �L�\�}�s$&L�YNw�_yj����&�|�+o���Qc��9Zq ��x)������8_���Rާ	��pf$�>!�����A��z�g1�U�m?� ���R]ZH���q�` �A��ʞ.�3G\4fû;�������G��j�WT�#�Kvɲ/*�tݫ]�.pH��S��@C��jϮ�z�`��z[�:�5U�&-�|+D�q�mz��8�j���ؒ.�S39�P�IK;�@�#~N�V$�7c��-�|t�&.���6��k���,PE�ɳSD���4�ʣu��WOω������T	>P7�ʶd߼ێu|�r4=�rL�n�����A�.�Ǌ��V�t�Aa7���v������u��Ϣ�۶78��Pƌ#0v8B��h�������\�kT�����iS�U�����-P�����F�&��8[h�d���9�C����� 8^V�-��E�JL�a���Ե����U�y�4A��C9VN�^r�G^L0�xR���t��,��(�V�ۢǫb��Y'�豐��c�f6F�E�6�e���[�~�C�"�-���t�(����q(��"R	�z
����������o�Բ�-����a&d�(��J�K9`}y\�lRkr7�X�������~��/����_##nE7#�.&A���U!�IWJB`vzH���.���>@鉭�b8�D��e�BjQ�a���.�iH�RR�6�ƎK7�h���e�[BQ��o�J�*'��ʩMf�����F��F���r�!���	������ŐF�5����N��͍ׅ�*��-�{˳3O7�����Ű��&�S��2-q�!���@�ߚM*�����=pi%���8ʰ���G�.>ΰ����Q��Ugaf���YǕ�?k�Ks��3+[ؑ������_�0�V���yw�=뙫���j�96�������M�f�\�s��Y^�M�u2�;�a���G�83Uq�^J��`^_�n�S�/*�#my��O�4N��,ltYS��jn��#ߧ���G�p]l���8�M-y	0�]؃�U��`�A#'WG�_٢A+�ٽ�AQ��B���l#�j,?���N��mO2���JL�:yIn����?�Sd��
��dHU����8�V��@Ѱ���cjdq��!ǫ������?=FGʶ}�ŗ�D=�t.kQ�h9�_*eқ�t�v�R��|�F��\�]r�d�JX�h4O�����	���Uj^!��<�G�\��j�0낯�	.�2��}Q}��BK1�j΁4X����G����睾�����NM8gޗy����La�R"��|�̿��,'J*���-�̺���H=�M����T�&B�ǏF�6�'��=�}7�!�S�!�H���Þƥ8�x� C�)�+H�4�C�&f�F��'ׇ��u�����1P�����P���y~�fB���-4=44�]r"��->F�N��ā;��̜K֘�7S�.<~��)��UM�rf=�z���8t��G�}�׽��y~�c���̚4��b���%���	��|73#�+,�s�����[�0��I�7���S�2C�p�v>o�������l��x��\2Z��4�x�������C�jp�
��?���淏��'K��UFU�_4/���<p	L��E�/����XM�X��;�d!>f�p�lZ}��x��e�y�d£���yč�_ȋ$�"����DG�)�L���*ۻ1b�>Pz4ۡ�l�s�����H�42��<C)d6��T���U,xgi������?��CV�\�S
�h؝��Zwf
<�*�Gr�!��X[��9+����ŭ�C��M�`N�Γ�%�2�����H���?$$�5��CYT���xM_��'��DP�3O�Q�~��V��
�&�2��4#^T��(��E9�����iś4��[�#��O��f�2f��)�Ql��%��o��
��,��KțPq�@[��\���Y��t._/�-�����Qy\�`��e:�j�>��q��޴���ɋ�dH�l�kH�y)d�o�J>&6G06�q��|  �qo}(/�ݳ�h9�z*�,*R�I�Q��
K�|���΃�of�ݦ�D��Y�J�k���f̷�X��&���qD4�k�� �u��M���n�f�\PY0��/5e�t����/P�%&ۡ���ޡ�jM�y迯�@hz���T?� ���Qc[��c�
�V�#���y�zmۆ�ASR�����4�9�s��uz��f�?g�^�*
g�[���u'Zc{vX��lXG37�K���-uq��vV�n�����m��<lEmy���-����כ��`eh@�s 4W�x�(�^G�z��{"�)3W�Fe���#�2E��7V�Ҵ��Y�|��֘��^�83��f	��goa��=M�"1��l�B������*��/���脄:�GG�"�0񊒊AE� )���rc��2��8�[�xfLO��i�o�C ��Ŏ!��T��#��C�E�鉭F�l"mK���n|��X��A�u�Q�����=鐃c�0L�8t����:��y�q~`�;��q��j�~��y�"�4�0Z�,X��r�ǈ9�[{5�&Fx�OH��,\����7b��7,'�@�v��������w�PTHI#ީ��m����c������q]�<�q"��H�}���cJ�-ٷ���RP�8����W�������36�E%�����xY������?����e7-��R`�W���TJ��:�à]�h8����yqc�:�A�R�=3�M`q1���u������ V����p��@�	K�$tG�� �M{sù�e�w;�		�6��~� d5M�ģ��4>�j
*M5����y�fa^ܑ�x���E�`��[7�6A�m�2:�3�I���R�63�p�ƣ���wm��B�&�۹�^l�h�̡���Vō(�ʗpQu��MI�%d[�����(iKY:-�K�u8�xG[���cYB��lu���(���6;	�C�['�Z��T���Ҁ�\l�*4?�Hr׳ �m�^����tm�����{�A%L5u畇l5~)
��t��Wh" ~l<>�"�j񏱍��Q�]�B��_� �&tFM�q�����b��[h��;�<�c��o�z����a�iN�p���jL�
���=�3���[�W�[o�����D�
����3�ә��L������d��:���N�g��������B?Y�^jRyDN�`O��GO�̆�	��U���$bQ�}�u.�/�S�	�(�m�������2��M��Ǩ
�*�n�V��8���ޔb4�q��\�V��10z9�UE+FQ�wY���hP�J�t M�':��6]Unw�=�U��������C�?ӧOv�̦���N���M$�v�]��ȣ��6�e��?�L�Ϛ|��%�(rm�Fq@�����Z��GiW١�����(��^�h�����#꒩W��ë����j��XK�c&���#9Y�ʾ�Ui���_4��w��*�On1i�U&?�7:pn�8�P��maG�JF�J��j�����\���P�\↜����\�+|�{5�atQvn�  ���ע��� �4���U�՛0�O�X�&��aLo����<*
�<K}�"߭ac怫�8_��1�᭒��[���jԖ�������~�Ե7E�k���%TG��ZA�-�t�Ջ�ڭ��7h�l��`�]_o�]w{2�y�^��}tZ�l�)|�C��%����t�g�����us}��5���a��1;��1C�P`(���!��[T����W���P4�9�X�2��[� �*A�9W��U��n̏����������O���ڊ*zL3n�u���;v2"hf�#Y������w���Ͻ>.�p=�w<sܠ�	Q)��g�X����>{��q=��vjS2�"GW�)�@Ն/��"Ooo��7k�m�5�g���t9��IKD��H�[����pb|�i-_�/-�*;J�M�˨��_������XT_ˉC�����Az�SW͏юD��چ���t+����Z���^4��l%��{�)t�؏�i��,�Ÿ��s>��\ruW:��V�zYW���[:�n|��f���1��3��#iG�����ŶE�,'2����)��'��4˘.�2�No�>ԬEPj%�EF���dPM�!$�/�jf]=P@r��(ю�_�YyN��5�ٴN�?�B��<��B�����oϦZ�P�E?��zWғ�:�Q���@'�����M�@	��Ś�g�{�8�)�2���������h6�f$��u�ה�� .�Z���tڒ@�C���>��l��|��9��v�>3sf�������*�c/�<�%J�i��6�F�@��Vu�@65�������;��~~��ԕ��0Y�z��k}NY�ʙ�����NT�9V�{���-���у1�,8���.�D����K�Kw���X�������$����d.���!�B��(���x+	F%����&lIW$U[+><>�������(��J�"����e���in̬�כ�;��-��z�u*���ZM�y�ɸ\�KA��@?����E8��{�}a�B#ɾ"��VYث��=�W_���qy��.��V��y���e�S�łAr�!%T��<Ck��کy_�ea�*)�XJ�����r�ĕ��S���E����XyOc��n��ke��"�㘧C����`גdѢ��oRF^��)��&����\E�OՆ���C"� 	UP�*8��tP���)0N��I�(Bk��ԇOtR��Y
�MO�2��~O�%�.�b��������z�^0��5��ߺ��w}=%r�#�<;hG����SI{�>^$���B�����K/��ZǺ��F����ĺ�����|�����P�Л뵫�n :��`�}�E=	N��i����_��<�����$1��<�d̐޻9Sǭ�%E��ܝ��$�R}j�!�����N]� M�h�]�m۶��l۶m۶m?e�˶���3�����7��"��6�=��fMÖß�ރ����x�?��W
�ӵ׈]<Z-�/�y��+�J��7O ]�����3]̍FPh��<4;)�_{�~�'A�*�_���&B���/z�4��] ���]-�^=[vOD㮽��[��v{�0J�\T�A�Kk�z;$�3�A��j�����*ڋ�w���_�g���f� +��)�C�/W�RG������Fk�4��6~	�l��Et��u
���8�n��S�X!~P$9-T#�é}�A)�@u��ĉ$쨉"�pc�<pжk&6�.#�R�w1�V�I/�b�����SC��p�Lt�i�������������-n����}[H�Ԛ�Us��+��os���{����W���,q��y����%<�!����P]+ؙ�"�,a��wJ�{7��}2crC�&�O��6U��_�\aKz�jI�w ��t��7�?>��9x&����F6 t�W���H͖ۙ�b\��+f�,��8�X���������W��lC`]4En6P���s����F�ʝn�9�
�4o+)�Ie\�st2����Z� ���7
y�yd��H)��J�yM�o��WԘ�-؏�ta�qY�3��``u�����S���~�\и���������,�8Ĭņ�Ƞ�$P��t
��(���\P�@��2(�P>0��W� �J��Y�D���� �i�r7��m�DoN�̩���)�ْ�7�����fky}���LD:��ގ��v3��A�aL0�IO��I�A_�`�K�������v��={�����4�˫v��)�[�pv6)�}��Źz�w繹�if��ʜ���m����rO,�\�p�[ǎP��Z���E��I�z��Q�8@�ł����_��\Ƨ�eŀ�9���)J��ѿZ4�
I��~3��O�����G�
w�B#���o����_�|O*���S'HL�w�m�1+�׹�&����	���J�f�<$�#�,d]}6�H�@%M�Q�3/	!��p�4��;�e���I�\�8>��[�n���$�R��P��J��D������J#X.Q�$�befyA_�pR:�,�횗a�d�G�X�t�%���4X�r����eu�ѹ%�#r�{3�Ւ�JE��g�OD c��T��a�T�k�k�2gH���D�F!r�81��X���E��%��,pn�lTI �\����Yq;���W�8�+*GAI���o�L	��>z����1��\�ydڱ���������&k&�'��HL��J�R�/�E�:����O�-�W�*��Rʊ~7��%'��*z�V̲�%���A��6�.]�&�i�7�wdѮ��M�����z��]OOj:���}̩'��&R�̀XP�iM%A��Ji&�@% 蠐�����`GG;5p�`�ܞ^��O4�F{v��U�,[p.��aM�G���`�O$Y��Q��d���8z�#��]&�:BW���s�m�	A�c�8���$wN:`]Ogl�l'afg����82�z�/^?�2��o��IE� ٸ٨K!�jt�8F�cF�j�[��ĖM���0�Rݤ���"��v��h�~�:ye�CSe�P��������eU2�RoP��,�J�X87wI�O=r'Mڽ�nA��鍗Rqz��2|g�#�e���W%Z������j�󿌖���]��Dd��k�E�T�G0� ����/�P`��h�����+m�Q�3v��m~vu�4��k�rBS>���E>|0��V�G�ohw&�.�@$EF[�o�E_K��AN�M����8��nRm6g��L>�&���[Qr�}��86��I�81�E��<�+a|���cM�t���.\xm���[��1�pŋ6��L��L�	�����Ӏq�3ƀ;�EM��S�R�Lƍ�e��=���}ŷe=�WU���i���9�_����32� ��w�3�S��U%�t�WZ�k���)Q�~��!.���bY�@�� o�b�t.3��m��&-\*>_��V��������Gp.��o���S��o|=:��iw����T�	�w��szX�n��>/���{/ :#��"=HE��FP2�r'}��V��MT/�s��Y	u��&�n�,�oMq���rɂ�+)��汮�A�����l�Plg/~2���jn�W��=�&���Hk�%VU0��� ���Hi�F'�F�d@�zf�G�OfS��k"��WbIt�X��h8B�<4��Ȇ�H���Ys�⻼X�S,-��g�Y�^��,��A-u�f�o���-����
3�><Y�d�M�rv�H��� �^d�=�p�T�<�7�� �H��R�5�WU]7 ���<�d:W7���m����wew�s�:���~>ՁK��cm�F|�Y�9b	�$������"���W/YQ�\rODsU-%7�V.H��V�����ݢ��=�]�:�w�Kl��Me-Dz�.�C����BU�D��9H�V�X>��Q/���6�*�����F/���n��$��H�l�XL>��=w	�~Ȍ6�A�ơ=e�Y��DBm;�4.�m�ǹ��[7�!�i�ߖ�nǫ1��=� �~��f\a�Y��뱑�-[q��y:]Z�B�@&��On㝁�b��V~��[�y���
�T�q��B�E���FRd@�7��V<"�\,���O�^2UN���V>��B��M,p��a�Ȃtb�|�r�^)���7h��%�&����ٸ�G�kaOkK��@���SZ�=Snބɳ���P�.����Q�\�cӮ�r���d��X�PL��g�Q�PK�OP�ɪ�JK���o$�]RS�d�K�]8��]?�rl�Oy�8gjҏ{W�X�iO�E�M%y��J	��D�@�$�Ii
OO�O�A���3xP/����5��謆l����f�+v-M�����!5"���^+nb�fG��a�SQPa
n�`#�&@5Ѓ#�\��cY�m͆�uF��x|��p�w���KOkE!U��t����TX�	�Me���y\>�����@J ��É�b���S��Þ~l�:z����X��9b��Y�ck0�,; N�a�7V�Vz�2�Ҫ�x,��}� 7�ᒻ��r��R��7�ÃfX�C�*�)-��Yh5;��Z?�+��X��i>>��r��H�0�ޯ�ΐ�������4O�'�M�*[R�J!�!P��ѹ�Q�I����V:>,>��-z�Mni¡SCe=�5�
Kh���W;��w�&f*�!Z�s����R���o������.&#s@c�\�u��Heޔ�쩌�k���u{Is����!���/���L�H��+:9���\���h��n ���)�9��S���YZ��r0밹��&̯�)%����ˆ�nh0���
����ņs^$��H#����E�4ǹLGO� ���`|3n���"F�T�\���]�,ѳ1%�ߠ�T� :��0��āpnB�����X��Й%#����$��J1�����Z����׏vq��4� ���_)P ��}�7��L��E���ĉW��lޠ�aC����d�iL����<�(v���0�T�|�y�����a����W��5|Y��v�W8��D�� �[|�em�,�TX�

��:g$��swXW%{�Nk�/�wNT���S�
��rq�0F��3f�f�uXZ����0�'ߚ,�ZG��a��3�ꊌe�KD�0�C8NѵG��'	�s�D���.� %�Y�%�3��K��r����w*������Km�����4����:���m�X�f�����]	�1�k)n#>Һ^uk'w��k�6�NԀA��K��}@��f�8��匮�_3݈���Gk#v��i!��-]����d]L��󔒔q�
��}���Aݼa�f�c�b���<0��OLY��ͺy`���ހ]1m;�Iү���M贃��Λ�s�\ �H�6����yM�~��Y�
O�c*�fx#&�V�	���_F.��V3�eH`���F��z��ր���"��IM�u�*0a��J�+�����k�t/�qJE�Õ�7祢�a]��[uEZT��~��Z�v��[���
DE�V	�Q?+T�\�D�^q�iH<F���2	 �bS��e��bI��R��� ���aD���^��"%�,řOGiG`0ƌD���3�&���0�'���`�'�cZ��Jr����@� �b����x��.͔��
�����I��A �)	��~m�=��DD�#��q!�.o"�����G�K�c@ݪ��7q`T�KMd��q��&w��u��e[�� ��E���q1�k�L�w�V屡+�p���%Z` p�~�bd����#p�L������'W���fo�TbN���qk��Z%<�XP;���{�15z��퓕K�wh��b.��/&`^�'Kf���a��s'eǜ�Z�11�.�����ۨds/рyd먾X�|�٩�ߓ{��8Ko[V[��1;�j��<7	�.���k r���b�"��Ρڮ�>Ӯ��6����1q7/P�y1Pk�W�$�?�g丬���
Q���j����.����E��eU�6���{)a3���Q`���_�ظ*'E���@Q�]�s��*����������h������|�ao���Dyz�ȳ�?\�?Q��u�?�u��1�;�n�>�Sq����{����Ӝ�j��uB~��/>��O}�(��nD�^u��S����
� ��;��K
���/x�Z��D" ��w���rA(�_�2S]BB}J�{����ac����?�'t�ѳ<(=w*1�@�O�q��?o�5�|7oK�w�
{m��͒]�.�A�3��u���9~��{ ���|X�l&��3�bX�xC�|�ȷ�����9�K�F)������z�:�ܝ���~��}_�֍�i����Eh�� �qC�V�ž٨r�c�ԩ��V�d6�
(c`L�%��ϋ(""�����h���nO~w� �)�z��a� uD��=�ED����.71�8���A�+L(��^AG�d��a�Jj�Ȟ�i���u�a�w_q��h5�SƸܟ��@��Bd���}8�%A�B�!�$��g�:�K�2p]��G���{:3��XYԽ��F7.�r�ЂN4����؁�oN�a`@0��t+���P��h�����g�y4M�MO�\�������,r�D ��Į
�l�*��Ä�lŃ�l4L���N̷coZ�f� mn�����à�w�����0��G�gL4�����V�!�2����i}7�p�8E?��wڽ�J?�/��B�l� WF�������H���(����4�Af�2�<m��t"p���:�~k�음�ė��<���xn���7�����d�l)pc)�}�����/�G�%$����`�}�'r�$7�Jt��߻���s\p����5�\�_���H�3)u(v�yhMv�Y��_��?q_���_pS�ud����م�w$�&P�������0��Љ��2����'���^�\D+ ���ow����}a��'�/aK���܂��w��������҅Y��o���c���Z��_����dv��+�{�;᷾�P�F`���-!4J�7M�����!�(�1��$�0�b0���z/ڔ{A�[d�	�p�޴��AP����d*�hI���E�A��b8:>�����wA׶v��ە9��5��k�#Y|P�ٿ��À�����B��d%�%c�Ѯ�Ys�����wz������#f\��N<Ey	Ms
�`�Y&��_l���s���� ��*�K+�
%�V[l!���9�:b��p��5��O-\]�z���K��=KN��O���I�[A�����J��ecR�K�U�o)om�-�����ߩٱ�sD9��_��v!�oà���bZ�vo��
O?�d*�����fJ�$w�~�o#�������B����Kk���(��M�����E�A*��0��jJ��kv#�7�P�:^\�i�R�L����@����3�<�k�C]@?$�	!/8ywS���+��4��V�+�zMQ��������G�!°q|=1�#*0үx�wD��;G�z�/H/o�D��q�/��[@@�wt��A��v	���(!;�������w����h�����)��@`u��q��;�0��T���A�דM���c�uvM@�'m !}1�<�/�ɺ�0O`+�=�Y<���v$��n����Y߃q:M�)ΦĞ�F������3g���.��/�)�J/�+vvj��m�Aؠ0�:b� ��qi)o��9��zؑJS��+Z>@@� #m���.#,<ي��������)�#�K��Z�<
�"�)��~p7��b�Q�'_�_������� }�5%ā[_�$	�%���=1�����!���G_�|���U�m"T��#�x�\+*bZ8� ~�j1GW�dv�z���n����2��e���4UmW�H3�IL�њ�ڭ�P����Q�_��o�!=��$ڎ�А(F�U�E�"mUD��?� ��G�b9!X��+���s�Ѹ�F���ɭ�._ "�����C�Wl�rSh�@hMk��)a���)�h@u�Mϯ[�7����Qѿ+�z��#�s�Q�q��ʅ/د׷�CI,;�ͳ\�0f�R�]h����"Q�w���8��w��������
�(O�#�<J\դъ����^I�0�����BN��:-�����ʽ�l`�@H�A�9��=h�X��;Hd\�FH�bP�BJ&1J�g
��	$	�)܌��a�i=�#��5Y%~��(@/dCOJ�z<x�4����z5I����i581z�|)�h��H(��ܦ&|:������)����\�2�͚�"`��s+V��쑈��]�1U͝�R��r2YF?�-��ʤzxw��6rfC"f����,&3���[é�Y��h��/9��Z[$�K;�CD��	f�۰3 h�@��-�<��0�.�W,K�gB��2�G���iuկ;ݜ˶g��%���*L?"7B�tf��a�Ld�q^
:��.������O�_���J��B�m���K4a&T_d����dHM���=I>~���p*�':�m1|~��+&E��-}d���R�ʍbu�;�K�㾹��J�p$ ?2��n(.���ʠ�,;<������̢p�������O�����D~�a�/��O��B�sҬ�pg��s�Wz7�迧����ψ���_Ѱ���k����)���͚&Q�y�X]�y˃������{w ��?d�q�U]*rJ��xB>ٻ{p�C��D�M��n��g��m�4(�B�����%�>:Ш0�p��j��h�/g��������Rͪ��f�/�8�ğV��W�L��6�i�;8{<�!�p<_��r��2����@�|����aj�=Cד�S�Q4�$1@�$��D��P�����`e�6��`��۪��'&F�� F�9JO��8��v�NͧN�
�@_�h�ZP���#N���'�~�]��>���ʍ>m�2�"�&����[I۱��M��&��y���)����7ݡ4 �t�����m��\�UА�����d����t���j���X���xV����98�k&���x���bo��;{�X���m���z�`Ϊ�:�RK���$�'d:�=����60m�Ī�J}���^l��5�p`?�Q�UPîE(3D?Hy���#��s�s�����|l��,�>B�F��rkv��?d��b���|a����1vPX+P�_a�`�������#u�p����	�y�mx(�hZ��L�0��
$�>bH��F>0�9#�;���B�{\�6�b�r3#q�Ø���iB���W�V{�k�×2�����*��������c����9��/��Ss�	����DL۬1Ps��fww"4�7I�CзC{H |oZ(�yc�����7�Pep>>l~�}p��PS��'4L����{y8�O�V-`���ǳT~�����ߜ/�� ��i��������w07��  �z�<�,�o�iq,N&�t*Y���8,%M;�TU.��c��9D�+�R�����-���Pf��ѡ�:rz������7��݇�� L�?����K~���r����5�y!�Ip�a���4d�5:o�jG��|���c�ۚ�rj�Э6��]�P{E�����9�+��-�:t���0�6~�V]�?����fv�XP�R�V�OUn۾��kb��[|���4e4}��Sv�B��f�c�B��۟t��`��&����L��t^9'���'-���,ګ�B_!����3�#��q.'V����{O�.4�@m��J���zQ�9bq�?���/}j�Z1!��,�c�T�1��¡�>V��T�u��"��x����s�˕����v�V���Fr�d�8}gh�?�@Oz0Sl�� �28�L��Y���,�-+�~'L��:"_#j��6�a��V��T�p0`����p�x[pc�� ���h��͎�$3�T����ݝ��7���~450���Ñ��%'��fb��F���>R7��&��|�s���()��C������XF��M�FC �H`�9�^;L�߉j_�`���n? �yّ��_�Tq�-]�vGaf��5�E����]�ߌ��������	>*+֫M*'�++�"�ɷ0CA��/�B:�;7>���d|2mC�@�ӥ�7����_K+8��������E�J����Bv� �X����;n��z��$������h��Ai`�ف��f[F���u��!��ӛ#�w��(���wB����i�{D�iyώ+x�ǿr��Q�����}2B�˕I��r���:i��l���bB�AC�E�)�ʎ�pw�ɑY��X9�/�3�əU���|���@!遢w�ȕ�R�i�'�8��ܔ���y����=D%(R*�rg%A6��ϕW�Y�ƫW��������M�T�.�<w�]�G�8�s���s������p�?�5o�m��<���<�]ktZ�߄����%������|V���������}>b@Ũ �Ή�1���h����]m��]�� ��0���J���/߮��఑�����䔈�����_d���Î���[��P�L����n�͏�ӣM��e�<w'8�L���`�eK���	�|���O'�\w$g���6��?�}q_��d����5ްR�kkj�# �/��p ��H��t�M�.��SZ��M�����aF%rEMQ]�)��J��z���I.��K��5������{�c���`����������i������R��BWN���iN<Ŭ���Q����O��7�B�Z]d'��͐�Y��&�����*�1��u�*8Dwi��E�
o���Fח6t������v�������kW���G\�[�2Մx�����38�"
۴��&���[�"����"�CIj./�sV�L��)8mz}��T��Ë>�\��e��
��?�!���x�N�B�*�|�8� 
|Op0v��KH�b_P�Uݽ�o�gR��l����%2��&��:��@ ��K�F� �����Vh�a~>�k�qd�h��ʎIA�t�ĵa�� r�M�u����F�.#Ŕ0�b	�ƫ-��G�`q�y��RuJ�M��h�E��I���� ��'gf}�\�����|����a������������s�q�ڭS�b�o5�Q�h5�ƵK4Q��G���~|2�7��fSҩ[r=�Υ�MJ��+`*9no�К�V�[m�[b\<'���	a�΀�Qh]��ʩY|^B���dfχ-�	v�g��j�p`5L�ȡ���i#)t7K�P�b��q�%�.l�ko�M�61/��p�����r�Ȇ�u=v�B�Չ<_�c`n�!�S��|�D�VQ�7��J��,�L�h�48�r�J3]��T��2�$�4��!}xB��s��o�EvK��E�q~�縆��u0WV�#���R��s��cv<���Xt9W��۩!]�_!�_����l	�kc~9
�7b��]e���ŁՈ:9x�x��֋�A��3��_��		�cϦ��
�啱�P�\�3T�V��K�`~�����~�Uz�D8K��nٺ�a�p@�BOU�yo��6UI8y⃄�4���P �2Q��L�.����ndY��~�
ʗ�k�p��\�Ռ�25ɋxW �b>_��w�";�+��˒�h�;���j��°�0��H����_���2�<�q3��d�-�y�u��VK���0�[��vQ�rRW��$q^���TP�`��7^3da���C�Ɂ%���������2a-�Ff�dі�ҴW�3Ī4T��J��l~t��i��Ce"t F[��B�Z�%N<@"�2k���ܞ��t�ne	�1��BOFf�:��;dU	���YK���a9]V�y��dA�/O&�o@�����AM䄒�If�onsv� �n�n���#��z�Fk��)��A�e%	��N���\���X�(|N|����&���]�[�.������,���Z ��+T�8�j��q��b����|Xf=\�Ų��X�Vl����g�Z}I�(�q��Vk!��U�7D�{]~���~�y� uVW�0��BI��]1]Ûp}�f\p�N�ur�8�ڌ�-�k����޾R
�XkIv�\�+�\��p#���� �"Tc7;"���~�� ��������d�0P����m�Nè�:���?�1��3W���Lr�La�G!a�,��!d�ј)��,<��a��F�f��G���#?��r��YC��y�����?|P#�j�f�Yid��F�B^���h�`�~����� w`⠡��(��Y��~0�hu�n��'��y�r���-j�>|����Ä^�X���Hj,`��Jj$n����n���i���a�z�i����q�e��^Q4���ߏw�u����^Mnm7�
E�U����*�`��޶㜔z���q]Y_��i��ЍN٥�������N�㸣�����6����X^�$���04�2;�H�x��2��5�9-"23,�)␧P/�4�i�7/�R�׶v��VU���p�%�>���J.�.�)��B��ܭ9���1`� E
���+��	�����3��O����v��ek���>��&��HIl8�K5q�K�9��ݯ6Y9�� �_�3��p��u:n֖z}ٰm*���xz���A�WR�0�KQT�]�ͪ,Rݠ:%�n@�sp��ND&P@����Ȫ��a��⮧?z���Ѽ޵<]X��:`ȯӌV�n��;_6p��+�1w~������e7'��~��0l+�{���q|�{�,6���b	�3Me�����"%K~��{���-e����Q��w8A������>B��k�G�b���ċ:.���G��o7�Q�^a�+ϗ�i1�[Kkk����Og�U�ZZ-��x�\�Ԯ���I1b��?9pg4��3�k�u/��ێ�����\
�W%^_O�l4�33�lE��[�
^#������ǿH��cf� ���xOwo+���5tԑ@y��Y�q����HH�� mR��a�N�c�H����#p4)�E�E���˄,��3�*'p����WH�"_i;$1|8�{�p�X��Q�@'��]S��<M�=��(�Oo
%i!x/��T#BZ䦌����{A>�k�*�܃���Y�kdz�b�g��Π��㚥�,D�2���*���*�>�\��W9Gl������J�1�p>Zu�c�k�گe��4���E���GI\��f��q�`�6�v@�^�(ɠ��8FҚ�M�S�����l#���+b��6����n�@M��eU���H�=���hx>c�KN�)��mZ*���{:���r�F]���R6������\>f'cko[5x�wDpJ�˹��琋O���]}�?��H�j���R�����f$)=����{+mE��kH}4�	ʩrVS�n1�#�k�ٿ�%�i��R�Sd��V��%-$Ͻ�҃�d4�̜��.9T+�A�:�W��
��Ho��x����-7B��M^�������BB���_����gV��қ5�n�U�E��1�T��D�$ ��*=��3���I��?�vm��>���`��Y< ��߬��҉	ϖ�i	�J]���1BhW��si�	n����5�QJ�{z�A�|��
N���W�s��*�A���6���$�|@"��j�ƸSX��E�is�:�gϊ͜Hc��&k{�?�	E��<JHy"�y G��T�e�t3V�QL�pȥ{���7�J��+�.�.�PY}��D�/�����{���8e�e�*�r�ҵ��NS���^U"��ִ����:�D-�N�A�(_�dbD�j%LՒ�:�\���L� G{���Rka��ˬ ,(��5'H��+�~}:��Pc�*b/�.y��_�x�'B����CB^�����s6zM�9M���v��S�h�+W1Q���g/s揁���|��I Dn[�����@� '���7K�GX���D�.��pg�Yv0H~y�"����P��HeG�.�ӜÃ��vC/����h%��BM������A?����1ȠKNz�Å����!` =�Y�i��sqҴ��ԋ�ۮ�1o^�$�A���^�l��#�ܸxF�K����A���O�� �@�y�HƸ$Y� 벉c�"��7�>h���.�+�Y�\u�or\�@��a 1f���5�cjW̞>>,w{� Ȱ�ǗږF�pY�׋��p����*}�n��OB�	�F��`FQQ�c@�,���kPO�R���]�&�swS���O�-�����/��k��g�n�U�]sb�sj�,�,�P�1[m����9[|)�r!7��Y���p�c]�c�+r"f=�)u僲��s�O46]>
J�W���)���u#�^bwDZ�� ]rOj�W�9�o��(9rʧ��*��R��luR
�:BsXTe��A����r"�C�ְʈ�D�(�x�yn>�C[����A+��& ���	�v�ɽ�u�'����.�4�1�8�k���Kp\<�E3ݙt\�@x~L�
�\��ܜ[ʒ�.z���t�
 ��b�d�[���|��maS�|.��� �\d!��*T�8�#5��]Ӝ��{urW_k6=P�����7~��6�-�tp�d/6�
XbY���_7^�w�W�g�"�Ώ�H�2q�������O`i���1/�.�ё ��a����q�^>��y��߃l�羆��<`�Q�k���"ʼ!�ѱ��Ty�f�2��[���ga�*�������(�j�����_���mmm+�߮���2�����F�;���Ԗ_�Ϧ�
Aw:Yu#c����9��5���{�U�=���`X�``
����}?W��Ea�:,,���-+ȟ#���I	�ܶ>8M*�-|bFFZ�W�'���>���_�+��/rm
V���@��x������P��Q$��ׇ�EȐ�����e���X�;٤��)�2�g�}��g�k%Ym=�b4u��Oz D7+y{?4��ۮC<n�����V�iH�������:*�*��p�Tj�,���C �Wh�)o��cs���a�b��g��ks7^,ypy� �%;�r�Rb�@if[<Oݎ�Nw�4�j�b�,s�2IX�C�zrei�ז�L���L¬^�g�Z������YII}æq��8��928;!���+l��G	ĝέޥ����dj���*s�#2g��l�֖�:�cQ>
�-^�����_~7J"�9�^�xŋ09G�5r).�TS�@�?�Y��w�q�E�36뙱�݌�&8�_F�ԩna-�b�ew�a�j[e��U*p�ZD�w�RJ�5ucf�p��u~IL����ϋi׀�'a�:���"a��c7Z&*����\ع��IXJI����@H��Ʒwt5�6*��1�6�Ќ�׶5"�#}�|]�W�Y����'�cs|ni���=b��H�
�x��/T��"Z\��*	����(o}.H*�Uo��TL^+�����oa�96&�1yO�����? ���ʅ�s}��� �P�}�����6�[�����Cm��G!A���B�)�P��j���DՈ%���K��A�>8�E�ŏ�h㱚jҕ$�#�H�Ot)n��GݷR������r����t���\��a��c.w�������{���|���VU5|��̴�h(	i~ށ+f��0s�A�?�
~���IK����ǲKyi3̆{���,#�Q���I
��w�����w�}���q�A��u7 {��>��;ju�ͭ����&γ�s�������29�	#;���k2��	#����*���n��u�e����@"p����
S$�f�����9N�;}�̟�:�l����&�{h�W������7M��b6�Fʿ��_�,��Y�Lr��C��ɤ�*qie��B�۷����G76�-r!ҍ��_Z]ϥ�y�1YL�	5��6'IGrj�UӎG|�q�Bg���j������?�o4�8#�SB�0�u|~W06b��`�^?��A֧;KH�����	$D��F b�\����?��/d�?P����6<#
� �4�&
��� ��ɭ�X	j���`�?��ʣ��(,п%%&/Z'l�� PK   ���XKm���[ � /   images/e677f489-379d-40e3-bb59-6fe87b8e7dd0.pngt|<�����P�dF��22RV�!BF�13J�>�|d��RV��q�d%Y���>d����>�^���~y�����������j�����0�򮒼&FQ���"�	�~7|:�"{W��|NY���vT�w��X����hk�o�w����������B����۸�?t��wp~�
'��]�ݕ����z	�`8��6�����G�.~�w����A�+���n\i*�SubJi��m)^�.�aaߘfq���M��7fŜo�ç���%����i��^	�H�*Z�2W�����ٓ�2�F}&|�.TT
ؕ� ����}�V{�Jf``��.�-C�)��Yń��1�����t��p��{9���Ө�'�����i���mƱaS��!_V�6�m���mk�_�g��u�����}�f0ms��ߥ2$k��Ա��飵�f
��ved�ʟ2���ffggo�7����^4S���ԥke���G������K(�7I���ٗH��_��'Y��O���s��=0��؏������Tc�4�����1��^v)fԀ��_����7J�����o㧋�Q�!ݸ+�Jf
���g%�~�_��p���Q�^�v���?�nx֜B�G�.� k;���}}@؋��Xjj��N��)�d�Ї�F.ܾ��,�7Qf.������ߛ��\l�rp��l��s��{����,U�7����Z��[[��n���S�U��Ov#�ٚ;Ma9�=�Z�S=44�p��n�)��������c��m%&�a|���rӑ���˗/�W99k�e:�<��W!�~�+%*�W�>��
����j�d�n�ܰ������+�Jx	���z���-9+�Un*e�}[y[�����]�/,,�*��]�]��; ���v����>�sߖ�r����ɓ�Y�Ќ�������CvvV�޿�w���;l������V��M����p�C�ԏ��0������5��o*���l��u���Si��D�����8Qy�-w_z\ӱsvݟ�}���n�g��Rn�җq����zC��W�%27���888�9sF@łL&4W'�񙞏�����{�%�E�ː�'ࢡ��335��K p$�*�ZM����7��~�����7��g_�@w>�쏭��P}6�s��d;�6�,p�.�:�d����^w�L"�	X��sa���Ƽ�˯{ǻ�̍^̯��gbb
��L����g�7�������z�p���ޫ�v,bǔ.��wZ\to�[>���JW���������=zd��``d�j�"Tq��ζ�$%%�� �r�߿o\Z��<YZz�%�x�?*)�-U=��� ��oW�ڎ�1ǋng`�\̀��仜����|�W"MO)Y4�?��Hd��n�t� 	A.T�ۆ���G��3�

K����&IAfk
���|r�\ꥁ�Z�6�������q�`���A���po�&N��Id=�w�v_WEE���4q�� �����T�Y���@�9.;���'I�#N����Ce���R�v�
S�~�G�1@��KMY �~�2<�&y��eִ@��v֊�qgZ���oc@�4
t�G���z�G+ڃ�4���S��D�;;;�7/����>7�����T;�&hoʛ����/�栉S@�=��Z-:�.0C�a��h6Q�ϥ��N�RzAA����L�l����	��[ G�oV��yS�j	F���CQ��}&�p�Eg)#�����#7l���#+���/�u%"N\M�뽔�U�CuY�x�iijp�L�տ��?|xv��2�2f@^��}�}t999��t�Z�4�_8��d����������?��}>���5e��ۘ uf �	JK�#HK�*g�x� ��Hs��z����GW���K��1��{�����VҚ��&����C�m	HJ�u{k��Ͼ��b;�{�$����w�V�e%%砽yr�o��}�\}����ߧ�HhKy�:j�%6'��� Y�21����R��l�w�ׯ_G�TA��C߀�L�2%{`�����`aJ�Ɔk5��m.��6����Ǔ���C���Z��8�i���nc��l===%8	Xf"E�M��͛���@���(a0���w1TDp�z��O���^�:�V^�{gg��@���8xs׏^��U���km-kk�r�d��|���Y����^�s-�PD^�50ϡ�C��i�<%--&�ث�	�g�����^k��]�-�|m�B~Q�C��V��� m%8l�;��s��˛ž�͹�e8ؐJ�@g�p�gkUQ��>�A��	��%E755A h4`hlm�-b7Lgnn�f��Z 4 a,�C"���FӜΈ+=�q�C�{������кdz��Q��|@Y-Ժ�'Gs1D���@[����F����h�@'r��[%`�h X�r�iJ����h�[@$W�q���Z����b�6�x~" ����P�e�®~w9��Y����5?Yi��@��P�R2��Z)HQ�rѭ��{��
�$������3� �����~����Ui�'g����Y��pQd���--�S="�}�2$�Z��y �t�Hu�J)���P����I_�z��6Ov�I���~�&�V�'ˇI��RR���vʮ��{�0�Q+r���]D�~�)+++�R_��1�5Aӗ/�\0UPn�C y}v�Lb�x<[��T:��{o����� ~ ����x��\]�+��ZG�W��$��/��SSknll�Y'�}��T�Ї���e�z�9�p�����?-�����P��\�[�p��p��O^C�3�(*K��������꽵���q�W"viiiOS)`�@�s��E�s�+�!U�d� ��׮]s��Ƌ�-hG�Ǝ��G�|A�w��ճ�r�҂ܢ"��;E6$�����,P1<�:p�f��r���Pȏ�ul�c	��p��s�|�+���p�e؜*�dh�J����o@�
�w��w���^ж�p�xћ7{V�n�'5uuݷ�P��{��nl���^\RR�?[��7K� �UV8�~!=�=����$�X�r�'��/g�+�����Q��e�f��a��r� ���S��9���Mren���*Z�A؂�#�/��������^�X/2؜@@zb�k?���J�JN��0�>������L�q��Q�;�zHt��U+r\�J=<E/�~X\\���ᐸqi� ���!�<����@Bv��|,�� �*���VX=VQQ�����I	���-���U�v������^��C��%�Ѐj;_s�ޒ}���{��'�n� 9H�4������%|���,�`|kk��Hު��]$��ckkk,���hL;Ѐ�- � ]ʡ4�藻O�H����l6\gt}��5m���N�J����!�{n�h8:��̔�5�PS���\�?| ��ejj4���˗�H>읷���\�m��vs��������fTAA�L�	��ö�6Aaaz�fff,n���Ŧ��T6���pv4�ʤ#ww�S�o�h�� �*�f�U �9 6?�h�$�HI� ���悘������i�����%��������n&f�C�d������lPwi�V.����E��E��`c�n������?v�w�����#H;�ΰ\� ��e�n���Z�"�1���M�!e�EB�s�B�v����ɇ�D0�L୘�+ ����44��xi��8&~T�]���k�N?�����F_�U��,��r~�G�!?�vN�`]'G�ATB���7px��HA~�z�	�^�&���Ps���!��2���}�@Ǭ=Yfdf����O�?����x�<�nj� �<���#�����f�fz���i�İ�T�B^��zj�*|����3��ِ�}��_�9��J#/o�� �v��9bbb �J���NN�PU8;� 0�ٲ��0S�=��Y�]��f����7����R���(�V�|bT�� &�i�͂�n��QO��.KAt�/,/GONNB��>Z�j�w��`�0! �ȂȄ�j�D�{��P�}�]�]L3��k1#�yb;vXL�XG�4���ZV0��B������ș���@�r��AF6��@�8s�`n͖�78 �3t҅����O\��==�~�������K��A�cE��h���6_��t8o����f���S����#���M�Uэ>�&%%}xR-]
��₞~�� �C�ׯJt�!4!et"+++!|x��%`&4G����. �c~��^~-�YrEGc�b!|��Y999@C�Ad��A��� gz�t���M����9y�Z��y̠;��J�q���K�佨�*���36�7{�8�9T_�-X�3�" �0e��} v$�'�_��&�3MOO���`��(��������J���Z�Ae�IbQ�k��st£�vJ�+�ea��l�fVj��fx��ƨ�P���l����UG ?!]��� �������2����$?���,�-(L3 ~A�.5�Ta0Ӏ�7� �1��t0i�L�8���	CH���/H���L�ޑ&�XAPR�AK	�YZE&��e����嘸Zͽ`����O]�'do���'�t���!j2���݇��aÁ�� ��в���=��GFX:%֣����^|�}���H��@˹NO*=600*؃?K,Ü���+����f2ek��h�)y��nCgﻀ� O_�����5n���8C��d�/)��M5���0α�~��l~|�����C�|4:���	{�Ook4�t��{G0�)]�CÌ�c�~kl��*�b9��^ו0B�~,p:�����?\��K�Fͽ�Z*�wָ��-��J%�"�xR倱��d: h����G�pe@�C�&��~�=�x����K��������1d0� ������:��u��X�����W7jD[�燶	�{�\6��8�������d����\w��h A���+ >���#t�$�]��_aF��&vo�0�R���-wq2� �<�QQ�hm��E�Jè��f0�����RRm@�A�����$���A+))��ח��
'��m{{>�����p���.T������g�`��9п��ŤW�>���R��8�
�.�B	����ġ�h �X_y&�0�����`l(�גޟ�ɗ�\:��&���,���;�����Z>{&��\�Ĕo'������f��n���Y����)�E�&`���rss� 	4($,�?��&��AS�����z�T�}�
3�^'��%G��_`p<�Z���g	
�\��A�,pQ����Ds�2
b��7)�Ϸy�1 �(g��nm��γι�F׹gsr�{�!§�lW����p��[�'�u�K�8�U�@�y�����#�̠� ��"��O���	��z�~=$Ų���.���`��N>���@֊��}���$ʗ�ѝ�ǅ��ݏ�.���H6�������&�@v�G���6���P>� $>R��+���$��.����k#�y�O�k��g���1f��߄=7&~����T��&>{��Z����ʁ�2m_!�T+�m�[k; � �Z�� 9W�\�Y����c'o[Gn���],[o ��O��\G���1|�c��7Qyf/���7`8T�K��H|��JC|����Sl�!�k�-Z-w�͠�@}n�1�`zkj\�V;��⢫�[��>��.=ƱrLW%����Ҩ�g���F>+����B۷E�TwLP6���������{���dX��QJV`> �͠('�L���=n� {�D�����,j<����`~��i|We%V�0���ĭT�Z���P:k^*!����m������R�������,'_ϥ����J������9���D�9Ch�e�d�:: ��d��5��<�D��!��j�������WK����֙d��"�pT��ᗉ���e<s�;
�-H�A ^��eŦ�w���hw����/�Z�*Ltt��p� +���t��{JP�7 �4�ϟ�j���2�W�`��z�a��w N��{x�Deh���Z����O�"b��]-!�?Wߎ6��7@��R��v&#z��������� g����E�����/�t8g�U6���CXo+��.�T"w�9����/�$��P�q�1���"XRt	6��j����;{U��a�ɖ�{��D
��&��%:M��=�#��M�9~_}�����lɶC�S�!P]���E�� ��L����X!iG���R-Y`P����&|c�Q��İ ��u���u2���!+��m�/�@�������sy��!RPB���Q���K����J����o#��9&�r3_l�vۊS���[��ց7��]fZ�` C���Mf�C;ހ���E�v�`V�����P��ZF~#!߽��
�kr��i��H�Z#(B�����,Rz=����0W��<���H��U�cP�X�kJ?�SE��j�ˣ7X������z�nVx;<^�vH�Wx�d(�s��f ���,�l=:�V��:��߉�艫7���@g��QԮ-(�7ݢޭ�P��𪤞�z@�s�~�b�O���M(�2��0��P-��`c�&��q��e*�災��-���_aa5�Ȧ6����}C�����}�}�H������1�";�b�*��,e��c%K�Ț���.�o�!�<k�5aȄ qx��w��񝳐z�v?��U-�-�#�#��/,u�	t�}9���ٲ�.��uӞ5��'j�.��:�Hn򣋊��|����8����1�Ac8M�Ώ[G�ʪ�ݠ1Pl��=�0��8�D7:�7���1�xs����<\v ��m	��4�U�(j�q\7H��Tr�7���֭��x�� ��.3���q���@9W�F��dȾ���W�$OE�M�R��s���>Ǘ�kl���{�� ��v;-[��Ԙ^@��I�1Nw�U�\Y{�#2����z�$�{~YV�v�C۶K��v�� �6���I�Ns]�6%=���7�)\�����v�(���~����zu��P��'��@�� 
��V�0D�n25q�r�>�0���b�I�4� B'�sn	��������0�e�b��Ƅ���a��Rá#� 7�ٴ�A	[/�5���v2#����	���[^��s�k��)E��e��wt� @�kܼ\Q���6��^���4!:X�ز�^�����4 �CA%�j
�ց�z�Wen�b���XXe`_�NMl��a'����P�W�J��HY ���x��g ���KJ�& <���'�1Ju�����ϳ ��F�=��v����eu�}}}%�]m3ΐ%B_7#7]x �ƭ�)��Ɩ�2����W�����#�3_�J^�Qt(h�"|� �ϚPS�f�Ds~�D�� �TQj��轹t��m޸@94�R瘿��JAû�[���cӈ���@�H�� }�o�pq�4h��������˪p"���'�W�G7����F��աd�j �WHf-�~��V���S�kY�8��p�]�L�f��Ih�w�%��}E�-�"0�t��m����^���t��K�F��*����.㷱��QT܀��g���D	tijB��`U�c�ѭ5�Ni�A�5X���^ph�A>�s���Ň�b�@ޅ��q���&uw��~%5A�P 6�9	��.���FI2�.�L���g67�:��SVY%'߹r�ޠǨ�ac�f6x5�8S���^gL#�̎� Px���求�	�5��	Ze�%�>�l�%{��f%�[�$"́��̐�h���+:�m8O���O�6f�^L+����cHqk����o3M)�*�e��mP����s�ք���f~���MB~�����!�t0������k�U��:��~�w��S4(�|e�9�����G!�����6��l]L���y*f�+��!�{��������x���tñ��̾f-r����E}����Iw"v�����Ҙq�������=h�����'�@>�
�>��V�<_,�
?��)�Z�QEn��:�P�Ї)gkґی�H`���X��y�L�C��)ST����1o:�TQ�j�V�H[�q#mG��Ϙ�� 1A�Q+�>��oA�Ē���&U�O�d�^�|h���(���kM��E�6���sW�Q,./�aZ7`�e�����4�d��L���Ґ!�_��.mLw�]�T�|��;������7�Sm�&��t����~�Ո��@�.�z�ih��~�l)׊�U����rA���;�`����Î��;S�jF�	ﺡ��Bd��b����Zk5�LZ.�p�x�0�ӓu����2�z���n��G+�S��˝�tív#~Ўr�'E�.�89'�,�*���e�@�ʃ�zǙ��1f��@���Z���}�r����ڝ���2��j�\�o
�'Īw!s+����cz���`���ɘU���2�zQ��G��r1��)��Ke9�A�k�2�������J�V;�F������Q����(���fM���.H���3WOj�'�]/�V�Ҫf�����f�7h�=1�٥G�������6�������X���q�f�Xk�e ���bʛ�^�h�(��f}��ȋ��"ۤ�L9�(��� ���ɇ�@���r����i�BE���
�5h�?2����k¹�w@-�,�j�+�^/���N���
u��p�DZ���D}�a��%M�{�j�0Rs��HU���������Zr݅����ӱ�۱�cO<g���A.[��jĝo�z��N�fP�j�oQ�nH����ɢբT�dT�Dro�TS�0�l{�*g�2CY#�{�*&�f�
&�n��>�-0!��D��.h	���L4v1��&�m���x�e�iOB�M���v?���/	5O-nL�
u���2^����t^ut]\|F�l.D1��Bg%_g���z�����l�I���P-9R���M&{w�?<�[SS#(:�*xt]J�����X4v�M��}�M�ۘ��>��̊t�����)��$�IT�Bk6�#@W�t�R�p���X��_΄�1��8,�P�)��Ȳ_��ŝ�U�ۿ�vU�� ��3�iX�y��s�K�$ m��O��~K͛!���7H�5�3�}s3�nU�:7~�?�"�B]�� T���mbX�4}d�`������|�v�
ؠz1Ѐ���W0E�M�d+��{��R�zߞw�����7�:%�ޏ�J��
�^��/R41�J���i�w��y0�#h�h*����jNR*=2W���+�vB��$*�	�n��m�{�E�ᕨ����H���B����Ё�QG> qٓm^V����|J��o⛳>��J�-�U@��af� ���V�-=ɖ��2⁊����0a����UH�)h�&����-R6ɲ�g��-X�6t���G��hd��(�'�{����:B�H���w}�y�d�|)��:�o&;��^��|��U�Z���)�3�'NR���&�_��V,7/B�xNi�aߩ�>���<W+�U�Șߢ)p@��ͅ�q}�z���IFu!��o5m���>�5�����=����Hi#Vn��.���Tgz��U�ҍ�>Y@�̦�KQ��k�ҽ���#Z-��%X���`1G��+T_��O�X?�܄}���n�W�B�}j�E?GI���P���}&��7�:m��_�%#��= �^������?.߿�����>ʎ3p����u0�h�����R�흸,�c=D �ޮ��٢�O������_KK}���ˮQ����՞.ǅZ�TJ$��6��C5���l�H���@5	��L�ͦ��'B�Z*��y��$!Hu�(ްq�da��
�X�.l��\]�~�
��d�X��[n
܊��^���@�����>=�h2;���J��g��0�&��.\�îI����?qBe�?�<� �ɘ�����b��,�����.���׀AeFF�lt��#�D}a���2)�NI �T�,�%�{�"��.�k�
�=
#^�.��W�G{�$~�]/ ���9�d`�n����#q�=���[�pӧf�,/}�����d_�o>~�͊8ć�vyrd��0{���a'�l�E홻��[ҧ���'%��9M�X�U��	�YL��0��/Bt����4��*�79�3&0����s�[�?���D������:���P��
t��'�@���
���AO[u%��A[�= �f�䄡2�[ ��p?��@�Go���`��`y��H���;�O���q��vrr�b�׫�j*!M@���6`27j�>��V��Q� ii6����Pv��,t�s��T�6zv��d̪��~M�����c�%bؤ����UL"�}�hm��7ڕcu��24@��?�C�-�������S�/�^�úΎ475��U�^��C7
&���:��E����(���|�}��~���R�/��u�Su�_���rn�	���$�(�1~.��}���ҧB��n�t����MQ��B��:(�}aU��,�a>~v��[~��~�y�������b��+3U�,�\���J��D��;��NU\9*��	4�#�!e�B+��֊y�x�)�u�P��Ex��/�A�n�tKl��n�pg����L���)>9MG�*����E����+��Gۆ�)�z���P���~e��`@|�=@m؃/C�I�ϫ���mnm�6¸xRZ�BON�?�1CO2X���'���n(�&%cY���{���x8+tUA�g�eA"{�Уv�Ŝ�Rb�f��(((l�A�
ég�X�Ⱥ��� =��g�И�H��#�Kq�fճq@.���L�������6��	�~׽�5��*6H�2=H�gf� u��c_�Wq�BF*9�Z
u��2d�d��_�{"�赫@Wuёl�p���e�f��o������������-^j+���o �>D3�C$׏P����%-$�F:�s���
"��F�A�ݩ��F�Ao+�*H�~0v_��8os��A�-M�f\*�kQ�8ʨ�~�B5���)�`��WV=v��������@+����:0����꩗c�����B�^�AF-�2G6��tτ�ڱm���8��
�Ȳ����
]n�;�
F��"�vu���TJ�@�r��P��g�!0`BOAl�����P%X��9x_?��Z�J����C��2T�6l�g��⢑@_���f�9��u0b��lŘ����	�`@���o��y=((Ⱥ��S	�&'i�h�w�� ����8F�œ` B\�}�`&l��C%:o�h�:�8�����?J��~R�������E:I�*����k�g�H�0[$�fg���̭N6 _AF�|�qv���q�����z-a��y��ۯۏ@8���J,����va�|rA�~�T��r bz���Q�N�P��.���N��͓�o$K���~/
Z�+a�3]����]U�����U� ɂ`}MNN�]����ʛǄl;��\(����_�َ[�żSmp �1"���g��Z����0��2:|ʽ�����G���آ�g�@��(�&	e���|9�繪j?���ve���[��qϋ� ��k{9A�6g�/�랣�cN���[��$]��rRX@Xf�V\AAA��86@e�M��	�R��k���0ϲ%�*��]2"D
�"	��,dA�J���1�>b��r�َA�@��#Y����V���&��mvIj�x%|����W�EY����^2��u���� Zs�^UK�A�@��_B���na���a�-S����6g���Tg���������5]_%a][����&~~~�-[�ܧߺAܼ�<��
P9��V]>���s�0�������Z.z��0�
۔b������2G[��3����t�%�U��7����Ub�+G1�U�����Cb���ϒB�H#����tt���N�u�_�4ܛ#K�~�"��P6@5��B��?8Z�,H�G�?9���P�I]�xI�R�W��/�9�Cj?���R'Z8"�EW.��f���$��K��]x�roa��(�]MǺ�_�|I��}����g��G��_ � jHKSK�	*8�E+;���l��0�7C�1O���b;lLo �����Jl�*f#(�N�� ي|1A���I�;h�5St˭�}b�T����i�s �
��Wf*����\gFe�̊d@0n#�f$(қ�P#T���6���ԭ�z�s+8\��9+)��cX%���C���	��f�����*l�[�:6P:��Q/��*��ά���Jx�AK݅���"�I)��OQ�-���L�O91?6�y��\����Yv�hI�\����X�֡� =g�k��!�����P���i����J��������᥎�Evs,`�����?�\�Z�>���/��X����'' �ݔO�ۙ�^L�Yk�������=��	�6OS�\����}F�w�%�A%o䖤���Ӏ*>��ݡI`��?B�,� �l	��>^QA����elO�]�ʯ�|J����sMSA����A�s���/���M~���OuGĿ�w���Pux�ą��]k����)b�f*1�w��h�#Nލ�ۢ�XL#�E"��r�u��cs}��Ņ�';v��rN��,)vk��s�Fr�3�(�3���!QD[� �����މrB�����R�2�[gihh�Ƣ8��B/����d��\!��t�>KŴ��[�N�`�vp�>�i�ޫ�T�rՍ_�!�7�X��|�#�=�r˽.8ᗮwo��V'�A�Z�sh�i@���ǜO�>u�n�����jFn��A3<2���<5e6�utYF���썛��G�$#�~�V��n��4(�.������59H�Ѱ(���}%��>7�("������ޙ�qN�hk/	�
�K7�����������̌��G#�x����"�I:��_�*�%7!4�O��>sP'*0�Ͽő6��e ?�?�f�����|(��q���<�h`B�I��D(�dĸ�ɓ(��(�i�\�G�H���_�x!Ó����m	���vzC��M�i<b�W���8W�k7�j����n��zqG��k�Rv�J�K�\��Ml��=��l�I�
�����8%���h�{Wiυ�����m!{yHĄ���r����)Y|#1�(�5:��鞐���>4��ŕS��i���c|�l����ߞ���w@b�ӥ~��/"�<�D�vlNk-s�`�,��(ߜ��>?JFC�tt�6ZA�����Ƅ�+�ǡ��~��O����'7�X|NGe��-mB�&$'gefQRR:b�%#���\�T��}sV��?�<���(BWq��&�[��[�ð����<�c�&�>}��z���V�
��l��,� ���!��Ҭ�rh����d%X[666:��ʄ���ZH���!�[X�`d�@�������?ES�B�ԯi?hj/�����W�A5� �1� �r�F!�hL�Z%2Y_x���C@�cӔ��{(+\��i��@?6�	��|@ \e���?�����=8x
�gbҲ��dW�!!$���V��]z=������bs�ܼ<Y}��K��k�)��D�uW�v�n�td�s�YZsl�
�����_&b��Nk/|�̯dHU��.��n#�$���Ӓ'a����İ���	�9��԰��#ݠ8~�zU�ea�GGG�Ci�?�q����O����^�ޖ�Oȧ��3�O�d@�0�����I�J�N���)l������q���^)4�waJ}�0�+Ѽ�;ѱGΠ۠��k�S��T��f���*��^AZ_���>#�bXb�Q�=O2�E>�2+�5
5�)1N~W��׵kr`�����J(�Ql/��q�X�v��իWϫ8��y$H��"I}<>��8U(�;Ɨ�����̕v
����|B�a��k�m�|G����͗�KS�8��{<���?�2(XIF��>��E���3_ ~��(׿oV^�o�5x"�'&/�6�(��+dV��L�������W�M�g�i�C�Z
|���y�OW;��ƶL���o���X�_����v�;����� ϔ���4	���,��D��^�U����g���5i�m�����3Ϫu�B��5U�vX	}~4D�_���[�aK��e�cO��T�������e��yE�z6��)��K�hx�_�s �Q ���%��&y�q�"��Y#\I�	�J\��֟�̺:������k���:�Q��3+��t(�u����r�&:N���r��������_�rV��C�Ӟ�<;�j��ϩ�{�0�3؏ԉBG�%A�@K�_��5�S:���ɾ}����($j�g�,���J�k(�@�1�����ǋ�N�+*��J
�e����z��2S�k�!�=Wa��YaP���  �sL̟�Z9�Nu�"A�K"saU���Ɠ!�C!��o�`�P"d,-��y�nA�m%ꄟ�3dw�*���������Y�Xi~Lt��ؖ8�l��8��/�3D>tq�m�8�t�ۊ.N�bv+���VM�Y��jm�����	FV�xG�ݝ*�y.;;�dD�$�S��DZ�Z*"1~v$���ɱ�ȯN�qg�֘7u�����s��<׮Y�k��WUU���������
m �Wp3Ap��Iȵ�,�od�����|�G١ZU��0��{�][�
��32JĒ�5UU)JY��%��z�1����R��֓E�0ѥz��ee�uu&���H1X*6  ss�?�x��qp����_U�=���YAl�5J�H\�$nש�At�������:@�Qx��#5��%Um,p�j��ȏ_[�ry�5~~--Z�y��݅��ɵ�p�y�x����t�7^v�v�HF�����`P� ����o�:��%#]����VB�샩�͊6��h7F�� �b�%KLL,���7�muuj�Y�$��zz�{(\�j%u�	}��8 ���u��@O�O:�j���0d�u�����OX�YqFA��;K)E�H*����L@U�;�L���ڍ+��I����i4+o՘xĽyt-�7�����EyF�a��!�ڕ�W銵���q� �jc�����d����:���*.�p��:/��9yG@��41&Ϟ��X�u��/u}��o���Y�r���^u^1����x�F�8���%�6Yܨ_���^� ��ر�6�g�n�M�[�f;\��1Di��{*�7�-�DL�>�� ~Bh+�������ʇ��Z��9PV^�`+�f/'�s#:-,FM��5h����M�G,���Z��{�X5� Ԍ=�B;Tdi-�������%׾���7��m
���Rx���xTms�kv����-�qXR��?��S�7~�������) �b(XMf)����<����J�>-�e� �ݲ�6fni�;�zE�E��b"��(77�k�u��"m3f_�����Ȅ<e��0%�?�� � ���ڎO���Su���;�ig.>��GY��L�ك�f��Hm
r1�_��W/\0��T(�Ǧz�ѷ��	Y��e�QR�����İyKL�=G\�i^ϐ�PV�����Ȉ����+J�o'@s��|U�(��W�Ͽ�&�}��$��^L���\4^�x�X,���s��Z��׹�)0�Y3V��ܱ�Ir�K.�� D�o�x�7z�gt�S�Ja�<��Q����.���Yc����!��0��?}������6&{�ѨV����5��0,��谀7�/"o!x��P6���?a�ph���lr���Z>d��8`�JXo�����%��BҺ�UU�tg9?��Á!a�v���޳�1��>C�
O�� ���)���PV�N5�Ӗ\���i��\q�++-u�a��u����5�4�ǈ�S�A�.�!ڒ���P������§P;>=k_����+��#?�����/��pq)d�^�e�n:�N�]� �������/J< m:�zvmx��IHdu-b����A�� P�tu��|,mr�HJJ��'/^m\���V�(���|�,���;{f����i{��'���2��)�D����ֈ���.�y���<z��f��V$ ��ōpm���˥������E;n$��VYooL����r
F����O�Z�	�6�}�㕵A��			���Z�SSUU�����s%��o�\���US*��	q�]4���̇n4q	0j.*J�������[�AK�t�a�QZ؜.�㸜s��òw�J�{lO�N�"��Ă�a9=�sz�!H��y�=����[�>@�>�D����������@5��J�,��=���Z�4����TX��VD-)&��H�Z�[��(�;��C��j�����y����]������������a��tP�'>�#��훁ֱ,���0��QZ��T`q�����Ǒ�/�cw�T��W�$
�^� ��[jY1Y�m�nZ��,�t����9i^��c�;�ml���l�Q�o7��~�V䈐�шy~kY�쩋�#Q�t��!d�r�ɖ�ŀ�Z�'��������1��[gO�zy1GFF~������փ�n�d��B�>:N� ��}�>�ې��s�۲i8G�Յ���������Լ����^�եv.��g0�]��(k���kz?|Hd,��zHM�ﶶ6�_$͝�F�rdY��2;a�����˗D0P��[�&�� !5Z�k �^"�m�M` ���V�������!*���TJ�_�pg�l*L�$3E+ t�>x���.PM����]/j�����{\s캒��v�O�GQo,�cM���������l [&Nnm�~�4{0{�����^Э�(�8\�>����Q\���6��
�����7�= #:��5ى����Mrj��fY�q/{��y�m�35��"`���gc�vsW'��WZfڒ3�������)��⺭�<���56����!�e�JC�x��K.�KN�V5������]�Y�J�U��J'Ѵ��>{�I+JUFF��޻����=U�00��D�oS
��Nۘ��Ά�^f�u��=+�dMo ��������b�ʄ''?,˼͙^�?m\�{�����u�0�O8W������	��������zFF0�0-ON>tuu=�\o_��F���ʒ]<G�V��rO]}�Xl��x�Q̢����㺔?��/o������W>Ps,���2	�\��k��($�3��[��DE5�)���SRRn���^� ��;�:&�
�wY�ӧ����y<�B��C!�����䍋���W^&t��4;D��
�'�(�fd��
��`BKK��7�'��|��<R22|��n�)���"�q�{���[��O�Lk�j�f`���T�-Gܧ�V߼5��k\�_T�S৯�`���`$��|��˞�����}U��n7���K�˃�>*ٚ_��}��2�����FZZZzH�19�����asf�L~��l����ܯ9"RI���]Ns��8��E���x���f�Dv��s,���
����c.n�8,96��5���zy����R�f��^�ab"Pm	����ӄ��%	0�mwx˭垪Ɖ��~��u��,U<�%�]F�~?Wo�Z�ܡO
�*{��~��F�q�1�CZ�a�m���dـq<��
�.���\g�@��XR��!�A�'�ݨ��@��d�Vb|ϯ.�j'/;�D�`��b�d3�������h���]-vg�u0���+���?����n{�A$��F�C�E�iA���C��������f��R�\x��>�}�r�{�9�x���9��f����ϢAX��r�w{��;aW}lgL`�.Ilj��.z՚�2��>�uWp$Fl��Ԥ��d��G�'x:�
���#[#&~ ���$�>|�0�BFF�=;��^������;e�c�3M* �/��.Kf�JFgffn�������Z?F|P�4,��k����~�=[��P`t�൏N�N˹�P�׭����I���>��z\�9�P{[�`�����W�|4�|���Dp�g���DDDn�ME�2
����
(�����:��bl���k���%ib�IH�T��^S �O�5fv8x�A0�t��OÀ�XF������fVD��G9�,,�ńhHi���=h�d4������X�1���fim}�llj�v�}g�2��ގ�W��������X�#���d ��MQ?�7W�39T�
�_��(���W������	�	p=�l��W-wW�d�f��m8r���jͱAAE�:�l{�!77�ֆ����'xXߖ}f~��3�}ݱa��9{�_��ׇ+�ˇ��j_BXW�~#��Jθ�
B�����f4�
�}ɷ�WnJXF��9�܉Ҋ;��=��CK^��H��OB;9�(�hk�nf���Dº2�cZR�Ą�$��"*g��=�J$����jC�l�Msϵg?20nes{�fd��n��d���|ˀ���ᡔJ	�T��S�>�]t�﯐�8����$�ۆ��I�#p��af�oS�q�ё���>��a��m3������҇�M�fy���������u,�9V6tu����>*M��"�5�5{ssx{�/A��C)��ɬ,�z3�ĩ|����+�B;}�]Yvޜ^��a8'���aP6c�{���e\�K1X�O f�<N��4W�����gK��\�݂�
��͎n��u��R��5M@@�=� �����dT1���!A�R ���*bg�><���י�{�I2��r���D�4T��̑ N=<<vM�B2m��9�bc�57�H�����d�@R��o�	Cqu[�������~��z��m�W�`7>��,�:f^�=��q,bT+Y�`rt�uw�S\cs�����j����l*K�V���>@q���X+Y�S���H�- ��s����wrz�$!�:d �7�@:f��a��_�qhih��ˣ3��T��À�� �#��gA�@²�[���\��NA�ۘp6����p}gH�|�ː��O����1�׈^�	^�kkk�w��;C/b/c��n��9�F��a�K1���'a���L���$�������(�,-�k�߈]AkZRR�����EEh ��JKK)��H/?-�����/�=\�@��것]b&���v�� ���1n�����������,O���_[-։�����]H�G�g��:��h�V�����m���ە��; s���u�QDkg���q�,`h_v��,"\~y�iZU%�%k�]Cj������A�v�歹�U@�r��������)ui�\�~`��'
��������9 .��� ��s5\�+]4��o���<��I�/*װ�X7@�N�G����S+Gߪ��
O
��SUSSPT���$^�%!!Q4+,(05;*֬)kn�h��|TC.,,��[k����l5�Ȭ�P��,��d��!~J�VR\,���2۶%DiG�R?6���G���XF�g`d
��}�hF�	�P���ޏ��ZZ_23) �0��=S<?Y��o_�מC�u���p~�|�80 ���Ի���䠟�����Wu�F{��ºR�_�d�Zp-_\!�����������'���_�����g�1<!��jk�e�p:;;mx����������������	��(�E����g����߂ݧ�������C�و����1�R�X����-���d���)]/�!�+�פ�� ��[n�s?��tv��OM�Y���2�{9c�����T��`$����.����v��B;�gg���U4 �n;C���;0�>���`a�C�K�͉1���Yr��v��~D| ����|�i^�C��� 9��U�PxD<d�%P�44P���'u����M�#�G��o�������2o��,��@���������!!��3��&��.�mt��� "u�X?��W�F����k~>e�kT�=Q^C#dtT�V�$u1!6�ըB�3]�j��\�{M�w<�]��>�/g�B�t'(�	�RL"��EE�%�jJo�$(f�a9 ����KiYY}GG��)��T�3^q��D��ټ�r���}�E���b���9�b$LT��0�=���a�0����`������_���/ד�<���7��_��]���'Z��OX ��΄c�d�&)�g��B�����7�����t�@G�jX2�Ut��䧺v���no8h�;ރ��`�B ��<���TWӸw��̡�ML$�p_@A9��\J�ZPP ��J�����fv"F�ȣ���	}U;����z�������Ȩ\ߧdl����w\�����+]a���s��=��"R�OH��X*�Ce`d�"���3��K��!�W�}}N7W�r�H�}��¨�� ���0�[R"�븧�]Hީ�?�ϙ�*?|�� �tC�L��+f Ƶ.� �i�QB4�U3�hA�m�6��x<4���X�~#-����G�3V�k�zN�c��g=�[:��F�Go6_���,.�νeѪ���8qrjai)s����X�����ک��Atr�0+e55���?>��V���X]�>$a�֛gg��؞WZ�022���	����9�,)��6����� N@bb�/KP7�>��vB�]�|'&�r~E`C����Z��[}l�X*H���0eG~���eddx��Ѱ����|@�7��4�ڴI�����nڧ�����u�g٦u�f�岗�<1�5k�6du��';�v1��������''��λ.{GG��8�^��n�G��
M�U�?yBhs���+Ի�I�Im�п*��q�����s��IJ��#a<Atܫ�xh�ϙ]�z]����LtYXБQ�6�g����Z�"J����rh�#y��<���t��,mwk�U�-:�v��VU�D��&p}m[����/_���?����
|i<��N��ں��x���)MfGŌ�(g�9�f�U��gd�7���ZY�bz��888�F��:/.x�����`_��,��V[KKKKK���^u0+0�)�?ޣ������1>�;�ҽ���0��f����e��{�k��G�d��Jy��|��y�W���>������u�mX_7�*�[xi�� k��@M|���?�/b�����8��6��G�]c>CF'D��J@��9��,�s��M�G&����g��䋠�0��fIC��+�:��!���͛�X��c��p��HV5�5�^�	�U��"�f�`�����Z��]��m�}MN���V�'UX�q��vzz�?�U���A�ؘ�j����E����9N���E]c/H���f�p9��2��H���-���)���I+uo%��^԰���7��?�;�z�23/oO�C]II6��E���Y;V�monJJJ���������xl������M
��W��oVO� ��H������J�A,k�n*��r����٩of��[�us}MS=�_��pa�J:�i4�dѶ�6Xsoo�L�X�LNFF��A�f%G��4��0��NBS3�r������=����cK'�@pS�f�+���ѷ\���ŖϯrƩ��UOU͡�P׭�-h�&�V�m�TԼ4WT衒{sMB1+��M��E�x����̌a���H����{Mq��E9�3/���?�yV�Nbբ����㲆WۧTJ����9E-�C�p�[Y�����Ydȫ\K��dw�P?�R�.q����¸��]L^D{��p�L@�Yz|jZ]M
�*�l�E o�'��Q��&�a}������ޜ��[N��Ni��d[���#���}߂PՎp��=?K'�����Y��Q�W�`�X@@�nf����� �h	}�ind7�b���t} � �uq�'�|Z'�8¥ϝh�P6#\900�y���l�����+|�:����J��ۓ�b�ѬZ�Հ��e�����Up3��0��L3�cBĞh���N̺Y��߬���}���0x�:�	��������T2��p���*�O�`a6v�̫Oj��l�ԞR/bz�#q6���l3��U%��3,/��"@�6l���I9V�8ɥC���Ϟ�Y頢��'926F�â���+2;�CDDT���������=R;8:���B#�.X�+55z8���L�j���T*bl����ԩ~�2b�[��������8_�D�jhh(��V���7V�jƴ������2�_�h�!<JG������vU`����A�X�'���(?�c8-;�j����}�IGfD�\Rؿ��\*9������p��&��"{| ����ϟ?a~��S1��xO�;�LLB"8v6q^El��v���QF����ً����s�;�CY�R�7ĥl��AӞ	R���]��̎�h��Ƶ�>H�Q@A���_wǿ=&'Q�l�ۨb�n#�o���FQQ�AY��ڶ��Jw��BN>�P ���v�r�d��'�Ǖ�J
P�	�R3f1��s��Z�&��g/�o����51��^���s`xO�n��
&D��3}tn�;�BYU�4�1����,����~�
�=�s�D�4����!gbp�"�Tpp�/V�,��s&���6䜉f�����9-0��Y��Du��	��7�PGk=��dN�
I�����.N�[Y�Kc[W۫�y+nR����41sG�К���\����L�)-U�J^O���Y]Y�����(Gw�d�}�]ǆ�n`�w�Q�?y�C�s$�9S�̭-S&ff�݋l___�[��U��u�M��LLL��ʨ ��:7[ҳ��sm� �^�7AWo@�5����	��Y���i a|<$�Y1�T�n���a����T��#y/5�����y򚚌q���//V"��(?V;��緁�r�lY��b��
(&��9��#M��! b�.�����n��-kEvҶ��A�\?G�oIikq�H�mIc8�<B�f�%	Z$.�^OT�y�w0�"��W�#�>���ui����N},�˧��S�A�y�X��I�f�@���I�4԰�ks�{�?t8���B���Oj�X^_�ƌn���Q$JKb�ɽ>B���'��8`�Q1$P8'D��L1����J���Xr�%$�AMV��$_x��B�! v��)����Jd�K�e���z����K��Ͽ�*S�����])��}� xz��j��$zg�X�p���v#$�V��Zڞep��m���e�#ET��M� �h��}c�D�}�\ ��{�V���M!y�$-�8Y�oϵ}ǈ(Q�����#��ǱR(��������#��;��������c���'�ˀ�"aH
nzh���:��%�k�V}����3��~��� �qM��f� ������<Qe�GC-��{���B1�O�$Q���޸���Ǚ��ȅYM����1g�?:h:'}�/\�ڲ�j�;����F#,�����q��|*
ߢ�BPK��A�"�&`R��~AZ��	ހ����Q����(�^�xBK�t �&�'
�rZ�����s&Y�"^�y�"����;z�0�PYSc�'��5$pUT��̾6_g�].�}�)qhA��:��j?N
�,E�$������@�+�[��Du\:^:���|?#S,�)��`C3�&O�ǨV�Y
��F��y>^�J�r��]�"��\�f���e����pk��$ln��hrv�\��Ĝ~�gX��@�@�^y�B���F�:���6�ϛ�~.�	���*�{�����y��Vـ���)*)��� ���c�;a��fF�A��؄"U�4�?3��_����)�Hpv�x��GQA������X�����>V�ؖ��zb�ȗ����&�;��	��r#[Ǟf������zh}Y��藑+"�������.��j7r�b�>c�>¥i��D�ܼ�����Z�5Q6�\�����SMY��LQU����p9 �Pk<��[�ͬ��n�&%a�q��l����BBF������᭲N��X�Kȑ�����ίu�1���8�����
pG��˘9��r)<�Ue����auu��B뙚��f�
N��Wl||���A
r��MC}=�R�ס���d-��������@2��O��#�?r�LO-//��p��%LyEI������ї�Q�ի��`���g���G����27�td��9Js��$���n�E@��+��o�l7��Cអ����Ihrx���4t�7�qs{�a��D�ʸⳫ��F#`6b�������n���ut�>j����4��'��W�d�3<ȝ>D�����Nq�Ӥ�t↛7��JI�@AI)&f�z��%0���~��\D����[)��z^��A͚fd�y8�����r���}1ް��\_�-��C����ڍ!�흝���|2S�G9�Z0��/�M�(���a���C=ManT�(Ъ(�78G����d�!7�!��&bX"
��%��=�5m�E?���"y����v=UC\Q�8UYss8��T�#gb �Z���̵�z����C��Xf����v��ڹi������Qa'p��
��,��K{5\ykz~�z�I�'|�p�����	N03|��Z�k�SB| ��}��h ��":��Ry�' ����q�'��]:r���$����Ye>�79@�^Ⱥ}A���N��I���ˬ�G�C��nr&�3���"q�O�ɦ07::9q�b�b���Ց�Qt^	�.��V[W�.)�jh�к�27&��(*&���g,Km�d?�e�c�;tm��Y��ٞ��se�UV�b�����c��x�3M�O;�ŕ�Q���M�����}Z��.��~�vVT�P��˗/k�60�'&��}��ʻ�|���I�UVV��1#^EEE1mL.�u0����Ҭ����h����@�xk����͡����SA;���'G��OE �����<�|��H�9�D0u���b�����������|\�vMH��86x�%Jkv��(�l�6��w�$����ks��ё�f���P�I�K�1H<z��t�Y`@@�%����K2}���niրW�FM_��y�V�Ã_�%!v��הؗ�OAc�{�41=�d�<U%�)Nh�a����x�w���O��۫�;>�Ka
���A>||�V��2C�;$4JF�_^@��D�_�4�¡#L'^(3ĩF�lḄ�v����tP�|D����?��R�~�[VZ�[K%%e��ЧHa��99Ԑ�9;�?c��0�
j�=A��{�B<���	�T�r�_���z���z�$DfA�?��C�tzifVֻn��{^--�M=޶O�m���3dO�iJ�6jT�-((���%�������?�r�����jMޘ�9B��Kw�XH�9�a�`!����k�ߴN�[���8cxq��Z�ǘ�j����$
_���RuyX&ȫXU��K.��KN^I)���оw�*ߓG��e���~d�)����º��=*B�AЄg����=�%�~�ؾ礩��ө��J���$M%�B���6v��������aӁ&��I�Q�	5�[/=|����&���"����{5���V-���z��I_����k.}ջ���@e������ވ���ղQ�� �לA���h54a(���V����tą/������UJ�_U�����@h�\t��qr��)�?215�:��5ZxP$��mמ�b$����P����Pd����-}���k�8ހQ�Db��L 	>~���&���r�%h���@��G��`n/4�`,'U&LO;"��?f+��qFP`/�N銽&}��49$��I2���ŠS3����[ S����+�0��qqq�_H��R�>��x����� ȭ�)`�n���$@�+3��yh��-ų�����WΪ�_�<��V�435�29V^��u��'$80~g8@���,ٛ�JUMA��I��6��|�n��\�H�U`b�+5U�c�L�^KsSӑ�,I�h�ݡ�c�I�KPM|x���?p�c ��>��P� ջc��~75x���n�k����O+���F�0��O�ǧoUUUm�z��N�1�ߖ�
_~/)��>9<d[p?����{���t�}� ���C�0X�v�6M�ח���E]���w��*Niii���nhE�[?�3��5ċmx�vd����_E,��6�C�L��7��w�\b7�� ���ׄ�I(,ܰ��x�Io%��|�^�e|n����g�d��g�^�s'��T��k�쀎� F�o*�g�>3#�-��C�Q�U������/������Q;�@6�u\�>�|ft��(Tw)�v+�����㛗"��**��D�]aDBy�j��`�c#�����g��[���i�GB{|�A�jj����,�]��H��TQ�<ݙ�g�����߿ه{�yyy�&x�@a�G�D���O��x��wًg~I�0�ٴY8�.3�����y?����i�d3N��N�y|��.O�n���h	PNtuw�		����:A��^�5�p�N��"��6<���V�k�A�ronX�/���+pR+++�f��55j�K� f�҃�����m��o�����k�~��v�T�^mm�C�n6��o0������J�����&��U����-CSD=Q��Hu�r��QUU%�tr6g���J�Y[a��X��6�k����	$����^���_���E5�KR�T��#K����m���������������5�'Ph�hk͓����\bnA*����	�hb��@*����{_/Y��55�n`����>3�q���%��Xl.{��v���v>κ����#Z��m"Շdڄ�E!��u�#��qp_!Zl�i����:�q�՛7]%�AZ�;Q���*f,��"�S��M?dֆv����y����Ը3O.b�����+�.̑�9~�JpK����аB��n5���T��"�2+�uE'��(n�R�N6�Y��z}�:^M5�"��Œ'\qE�D����cYn˒T؏�|�7R�Cu���Hr~N�JCC����Կ������ȧ�t�oL �;i+uh��'�^�,�:C_���GXă�ޠh���n�!�/���@����]#�D�	�تR�����Ͱ֒�����""�oJ��P��ڟ~���@ɧl��͒����	���ؔ�w���s����>|����q���3:�q�
�\=�L�M��*�@Ӄ�t���� #[]QM8�5Ā;r��-g^�8��e=�h�3���ɚk�S`���Hʅ6�Q��w�(pQQJ������sͭ��|1!�и�ҭ�����V��0*suw���0�f��r��%����h�E����/ i���[��C�����x���Y�B}�ߦx�G8T�"H�B���̞#]H���c�?ί��M�Yr�i��*���=+�PSS{��EShÓrD���8��TP]��.пf�\���A�Ó(>x$߷ ?���='� %�O��ar�8���	� �ݪ%;;���#���2�Z�����+�J��:G��/�d��T� ����B,s�T��ۍ��""��\�X�W�l�e���% oL�;CÜa�:�
m��P�
����%J_U����E��H�=�Qr&��{��Q�p}b�C�s�U����/��������L�l�K�u�5<2�ag��,��6�>������x��S�[Uk�[aؾ��~�r}NQ�WQQ!�m0z}��khh��=<,;���d1��'��J-�11����@7���۟�$I�����Q��w���j}��C���ē�[ސRq猈ά�H�R��K:���3�0����-��mL&`J� W�3�JLB�g�ttTi���d�ǧ0D߶"�������yi�:S�+��F���Cv�e~����O	����(5����H �ͬ����W���u?lCV|����	�x�':�A��?ZwN�a����݁>��^������cu���XZU�Xp�:0(���O����Ķ
��t����-���@}��mm$�:Ob��a�������]��S�R�]?�;�8�p|0�0�7�B<�Q�dU[n�~�����*3KԻ���x�OC��BK�A"t/���2��`a��S�">�q��K�FKʙl��N����^���s �?��6FH��H��BCC�o/x��`��w�x�����*��;;;���  QGa�����5�"�~�9�������Ҵn�nd��2`o;8�88v�7@����Q��$oV��;��bL�m%>}���._����;�/1`����F��e����s�Qm\V�s�� �@5N��ﱤ�?f�� ��/N�/ޕ%��"y=�ʙ�p0q܎��I�^/�Ź�`g���P�mT��+I�h_���'(T�]�C������.ЃG��e��g-�>3���{|�����()�a� �Bd���{d�L�̠�k@�xd�D�%m��Oh9Z�s�.�
�� )M6�)}FRq�F���|�D"���T�.��V�S���ݝ����&��ށ���QE����z���'�ڼ�077wts�Ev�SC�� BZ��Xr��Ĥ����G��O��̐g��Suc#��"m����ϔ����{��(��4��+������Ν�:�7����$f���67��X���/���Y�� �ֈ� %r���a��	�~7�f2>+���V�?<u��dޕ~�#�i*Z`�bx�"off~1Vz�+C5��M�mC��ą+>�G��1�xި|�$�����M�K���G�G��jU1c��;�pqs���C�)~�Vl��:;��޵�1�e����-j���vX~>}���T	����㽫�;@�L9gz�LL�ot�o�̨CQZ����E�c�(��X�<����z�����nR7鄩;1-��g�t���.�0ڐɄ��ά���O��Dc�>������u=-�Ԁ�z�.�n����g�rh    ��Ud$���_%�Y��!�h���1zcf�������v@)?6r�p��_PӴ��؏,��'��7p?�3�T9�?f}ty�^C����l��������K�0���~_�>�)�ѵ?�z�g���	�#���g�B��2�Z�7�AWx����՟���x`�3ӹ��E�%pɅ���ąD	%��|ɘR	`R�\[��?ڷ�w��0Y_�X�YĘ%��~�%�J���:.(������gf{L^'�h�����	ی���xm�6وPo#ˇ���4�c�hp��_��٭�+D�spPq[)G�e�E0�� �+!�U'*)-�QL�#
�/��l6��f����T���%JҀ��&$$0���yy�X̔�H�y��򨞽Ybgg_m��i1��4-�jc����k��^���7Ë�xZ�A2\�E�>{p̹� ��XX}<ɧ��[��@�dz��֢A=N�V�ֶL�;�n�n���%R�+�T�ev�6
���@ãߝ�C��A���pB�����8K���r�Q���4"��÷&IJJ��R;��;Xh��Ql��������d��RP�*?.���d;T�|�����g�(�-R���ѻ%%%�I�PU��ieSL4���i�$@��J:ⵥ&�Z��]|`D��ZI��H`W��Y���3cp�B[H/-�e�n���ب7D+����ɿ����V��%^}�j+(�Q��G}l\\�|ي,�<�)s4�K�_G+�����̟>}�������я@�z�/�,��/��(ٟW�b��R�o��^�����%��|<���d��8F�۰�����z'�5e8}`V	��B���_K<D SAǢ����i���P�4�T�׹*ԭ��$3�ٌ��R������UHII���1r�ױbϻ��{Wﾣ��C+���.=Q����3�Y,�����
����%RILίm+G��3���i�N�Z��e;*J�RS-%eAԍOL$F��Ʀ�3�HjX3G��ztL�����zV���]o@fo+(I���nXDm}��F���Hϸ���և�YA�K����f��kH�� �=ۛ�{�D^U�)6���W��=ߠ������f�
A�KN�VT��A:��4Q�4�*wWix����R�t~}�~yZ�5�/���3��Ύ�v ��H�s�ټ뫖��бY�2����N��+��כD<��j�sq�d�E��m���O��Ɖ�}���e�����������*��l��h-~��ʿY*�*U�ojtl,Ubb"�m�ܷ�:u2���[p��^i/	�755�<�c�	Y�a䲚7���*I8_j�cxړϐgn=[��>VUJ�ʪ��%��_�D�O��'7�X0�3k��x�F�k��V0}��2Z�Hr�EU60�fҮW����w��Y�/2���m�~U��7,!.��H�m����׷��[�b=_���vM��r-A%A���/��/_�OG�R�۟8�:�!<H?���{݊�k26E�̑k�B��Ɗ$�C]�-�E�M�U˯\����� ```�)?�����uv)-)��cחԅ��]�ɺK����%2�,,�FCi� 3��������vg*
��<�]��MGCG�Y���Zڴ�Z~3�A�ۑ���8��sv�^�ׁD=�A,�j�??�d��o}���)�����
Y�.����5��32ކ�����Ȱ�Czu}��U�10(�k��0���[�(��&��2�Er�O=�%��y����ƧXu[��4+�	 ����e��&鬄IJI��ʌ����+!)	"WBJ*��U?��$��|~��)��k�svuu�SX(�eNE�/�NP�333��^_~K�G�p�����ϯ��'��k�a�ϟ�J�����y!Y��%`���H�Jҁ�s�Lϗ}\E̋�]����a�5J�����CS��A-�����JWX̧������}�9�TpS�@�������)֘�B�jV�pEY߿����� �~�?�z�u�<f�����r9`��@mP���z����v{��0������.�W�ű�'��|�D#�򝪡�F�n�f�?�������� �KK���&�2�h����V����)S$�&I���]�������1��96hwE�����NL������'��\k�	<����oK".~҈�OB��骪�l�Z�d��m̍���#"_+��O������J^��	^�� �q�)�A��?۝�]� ���L�~_1��ntn������iE�VT>r�]^��>�ܕ���,n�Z��_�5s9ee���xy$��gpSˬ�$H=eձp-!��Jf�m�Ro���6�z.��y�O�������	8r�����,W��F(��8�ه5���&�9ݙb,���Ӥ�K+���������!��k��	ГAQ���lz>�{�6@��Б�\=�&KH��T��b��z��L���;B�E�����f�zu�8���m~�WH���b�R�<��o������h���>HN�&��@j���:�4��=ۆ�3�����j@=���]n>�B=㺹�����У��Tsff&:::�Js͋����-����Dtyc�'��D\t}���o���C�E�냊N��
��(��y�9�@�����D��Vn���\E[�U__?��R:\��w0���x~��6iU�.;��\M�9+J���u����ȓ���f�e9J��Pp�UL�LS��u��@��I}����![	\����<��Щ��Rd�(R��@�?��H.@�tUth�I�QȕN�d�UeR||z��;�D)�8���܍ �Q���r�Ew�-���y�5������!AV9��XP8�i���Rj>o:�y�r!"ŵ�@I���6`U8~�vq�+�H����۷��	 ��x�N8��	�'����]'�����IK����Tu�W_W1�D}�*���7��ii�'.a�M�p=1I�N+��`8�
�7$ ��&⣣����B&A����@L);��h�]By-�"���9���9.Ꙝ��a�7@���}|�6bt�?�%]X�x��D#�����T3����/H�Ս�>��_*kcx������;�M�� H�3a5���>q֪�����":/Qb ʱ��6��A 8����,;��� $�cY>���P�է�~�M�fCC5�Wa m74߽�{��^P��fU/>���I{�>S�D!���g�#3�OOO�n>�D=�=t��#����{�u`���Wt.$zJ*��^w�y��J������-��^���up�������Q�W��,	}�Cm�����r�19<��1�DA��mvo�P(�R��&,M�dm��~ C��k�f�� /;wN�҈��///s70��ݣi�cs��q"z(���t�j�窙��]�g:��NSõQ�����jS��0�����	\fi�)μ�c����4���A�>�א��6B���Js��/�<� L䂞a�;L@@��O�������l`H���K�w��B�Rԁ�5H���oD'����R�Ce'��pK�ʪFC�R|���і~%%,3uvyѻW�rV��+*�99U$����5k����(OO�cTE\����t�E���vDy_k�AEEE׃TT�\`����v�v�88k�yiѦc�ix� �o�ӹ�	��<��H�}�*��?NnԂj�f���n�|?���<�	&tw�d3�nPH���h�{����	"f�H5.�����Z�ܛCFH����/�-�&����X�nH�#d�֟+�n�]�3���Y&W.���J���q����<�X�J�%�J"(����u[uo�/-U����v~7%B�6�]�+���$\��* ���
ڨ�|K]j�+�~Q�%%�����β�Y�4�������������ջ����%[����7p�_�\�y�KǄ`�y��Ck�[�T��u>�Vޓohh(i{���-����d!�M)�]%�{?Z��!�f8{��B�0��%:F���3��+��ho_-Խ)�B�7Y�����P�M��բ'�������"�d���j����#���733C�����CJ�>��
xldjV7��2ƶ@�:�YDt�{�)""�kU��t�-(/��JB��bl���0�&%-�j��!$$�5 ����OH��Q�ܚ�S������y	.�E�QeQ��`�e�L���b%�:��h�;:V����ψ'�H�t���J���maa2�$|����2=����}�ϕeNn�F9&nY9������WF��S�d}���`,Э�ihhX��:P���R�i���b���j�&nu1x�H�W������
&'0�}���J�n
������R?8�k�٤�4":�̤�#Ā�v�ǽ�8��h�N���.z��s��[f�6+(hj� �P������A��H�E������AsG�P�_X�=m%��r��U�n"��؜�N"91
�ᐐ����[�0���N��;�7����#� (��관R��j4�B������x ���h@1�� ���ݹW\�uTTT�A��%���3۟��NI)�TV�	D�pdD}�i��j��^=\!11��x&Hk��w�	+����pD$#�TB�~@`t�/��uN���� ,MBw1�7i�رyxh�T];:�t,���ՃVq�ޱ ���J����h_d��5��zjj#p�zH�/7f�{B^�5c���r���'9�x˟�G�"��
Q}�c8��)�b�DD2}��4��s�ON��TSSSw�l���=?�4��y[�Ԥ������@�0�e��T�)8Q\���o����L����s�\]��=�4s��C$@�of6aak��@=�%�w񦰏���Evw!F�� ?����'�\c1Q���uh��*�c���� ��2<cъ�%il�����W��ٙN���SWk���e�)����,`��Q��+��z�J��%��Q#Yb/�H�5G@�*��k�?$��$�f��stU�DSK�nO$M���dd6���F)]B#�Au)�D��hӞW%�G���D��>V+��X�� )��adbR=A�cҨ�����U�	�Xl��PI��eҪ�����..����C��$#����l��g` ��w��e����J�.tBS����P(Mq"L?�sڏ��׏��Җ�a!!��J���_��cz>V���/��� �dz��.���4�Y�Z:�|wׂ���!)��?��捲�y���	������0C毀�2@�I((D�	�����at�(��gQ(��Z_B��uSU�h�ү��(����yDwVQ�`/Wdnf�-�{�'
צ|��#��7;�q�g��H@@��S��~�V����$�7�gg� >#�ޗ����׉����@2�6�����3�q����U��,ҿZJ��-��ػ���2�t��-�h0;�Y��ք
��@u�9����xBULN\|<ëE


��ќ܍v����z4���ڛA�&䲹=짹�L+r�u
�eOsY'�<��*���QI���L'���j������aL┄������,ب�v�g�(y�c�|��g�_�x�ui��Nt%��x�u�"�6~�{}s�=��l@� 
�f�Y4���󂟛�U�x��#O��)��o�ʧ�$id���4no��]D�E6��'%}��W�|ʜ_X���
'������3E�ۑ��d���,��H� X6�쩨�$F���#��Zڙm$�#�~��ѧ��a�}3�	 J6��2m]]]A��Dooo�zwWW/���I������4���_
���-//��1�[
Չ�(/��l�Y/����(x���ʮ�R�|�պ���#
Xz��"���<)0˕	� ���dk,У��:�����a�G��6�O�O�y��F���P�5h�FA`�#�E�^_FGF>���������u��ӟ�-���_�� �z I��q����\��0g[�A��k�����𛛛���z�ړGS�U�k�N��M  ��᠏q���rs�xפw���f�w(��o4�DF$�0-��@��������"��zr1�.:�<���"A@r�ru����!�9'���p������?��&p�a���00B�v&�%�Ζ:2��`E��pޭ�O������+ji1��,v�}�?�?/p_D�]�}s~a���8 �R5�+����d&5����V�#��-�u��|1�FFF�<��Η*��?\P� ��h~�^�l����g�:�����x~��va)�b�M������[�w������W-/�a��Uښ�⭋(��T$�b��qػ��(}��#:8M]]�^�2T�7�|;::g�6��J��^�[�i&7��ǳF�n��-��||2}c�""���O�(�_��r�|�Ҵ���U}����Q�;6!�(z �<7�u�22a���3�y����~`\^��tk��4����Jչ-��n��W\Z:��x#9MSK�f��OH�S�?��;����אJh*�D�2C�lBee��Y�Pf�*{;�R�	YY�!�ؾ��������?���9��q=���x<�� U��Τ��� �_�yQ|��[��n��E�ѩ��c����;G�E|����1
�O&'�	֍[S���-��^��K!ıOu�%32�mH������ֳ��zb�����|u�U�۴�C~�s�i�W��"\wR�!����$(Ŧi`z�CRC#���r:�6��N���B�Y��r�$$%�r[�P�:���!�*�Q�WE/�u].�)+��i.�I=IEe�I~�z� ����1X��B��������?g|����p;e��'��sss&��2�ߖ+��D�d��}�ly����/p��م�5��8�?f��۾۶�R� l�rE<�ll�Yu
o�R����1 �YK ��Ժpܟ��є����t3c��u�K}���*�����{��a;�ݳ*::�f�WĘ��#-�.�'����O�9A����lw�E�� ��tJ�o.2���?q,mܨ�̓-]�+�Ș��ce �����&���TV�2�LL>u=׳ kTVR��?t�	�����U�!��hyh���"�wN��M9����wz�7�L��9�Ӓ��]�w;ߦ*��V�S��d\����k��߽{G-fv�ȔSJ��?��/��	<�H&���Tʨ����>���^��dVp�ΰ�߼���==��q*���7J FS�w4]г�P���:��dc�����n���U������/��x��U��[����(����ۀs:!]��۫���~�wD��N�N�U�m�F��������[�h``�ֿ��MꉐeRaa�}8*����i���&$Piz����`+Q�C�؃z/H�
ե�$��>�9��=y�s&Q���~~!ψORF�/�;���<ʽ�kUe� `z�7g&��(@���&��F�߿�hHN�N|5�z���i#��z�l�2�I={�=��?��S=�E_R8�Uv��+"
0.�ŗ���~���a��M���� ?��[�� 8�X��/�����{�0T ���&�84��^?��OD��@H��T s���_?�bbb�:t����+i�������z���������d#W�
��i��}gvB�5���(��_������RH&��J|�t�o�U�2=�Y����ׯ�Y7��H���9o�+�K�ٗ);��IS�5o���S�v�X���3��������;���1e]���>-^�9�WQ��I��hMGHe�T��i��w*�**$Z����Ya. `<�e��}t�<�N��L��� �[�y���e�@u>>>�)�FY�oT"��߾���W�m�5�ݕr���1���%=F�o�5x�loo_Z�s�ō�:p�Lb��Sy��}���T�_2����>����������ֽ�� ;@<`������Jg��IX�\r��:gDIpE�۷oՙ�"Q� ���6�/_�T��e�����j�MN�s�Kҥ�,���Yxn�/��zF^<66V�.}���ȏ��T�pK_j)�# ���|��XK��?��'��r���"g��+k{ݗ�g�_/��6��#K�iii���g Q�XX\b�a�7}�ŕEթ��OR����ozzt�M!@�O��K�B@P���Z�-�;q���$�ɫ�.��Uq_32�7� ���H��Vҷ��'��������`���H�?c�O �|n�W�k{H&^�z��E��_.JD�u�걠5�ʳj�q&}�������L&11�`^�j��?nnn�/O�R�XZrj:G�Y�݇j�	��{���­�?-��(��x�]E�TXĝI�����IHH��Q" '3��ćP�PYS�>���֗F(~��߉	Ki)��EB���:��poH���Ib�W,��C��22>F^^���fmK*�r�-����.R
hk�4�J�Y��r�GV���q�Y�vAK&��{�j������.pp����m&��sڸ5�^{;���_����`tw�5�'��U?(\wGG�
#���L��*�#3kM��>�ؾ�c���Y���-�:LݭCD������=�{�%E���4�\s�:ݴ?R	��r�E=5�|��5�9�EP��6u����~�ͶE �?��������T�+�4�͛h {�*j?q[��5������BPgD�ʋ�p�?�Ro�@����яJWB��j����RvaS�bx0�YG�mRo�+ئ���H�J�+�,	���x���F���b��Q�͋��e��r����c�&�DsbbHL�Ϋ�����.�+�����_��8�B�,�1���I����Ǳ��E;��,��^P�Y�ʾ�\��P�s��!�,��F�[J�K���D��'�]])t��FF�֟�pq)��6�@N\�����w�`�R��Z�Lbb��v}%�o�0!�T���N�Q"����3/_��7040��� �p�s9N��_36���ʵ�u�mo]xs����"M�ć���+��U�.�,�F��-��~=,X��JsO�V�奕3�?���LDI��w�Ni+�q������K��Md�k���u�F�â֘�M�,��"��P'��� ��i�I�=[R��{`u������`��ش�o�X^
��/.1\T{?�RS[��ի;�����^Ն]�N\i���toA�G�v��������x�O=����5e�nljB�U[��:ZZ�<����C�ᒞg^<x� 6>xdQm��zff�͐;L��>�.��ߌ�u�--juMu޼9s�ȑƞ����@~�+��M5m������CAͿp�����gQK�4�"~��wK���Óe���9�:���2���y��*�-������l�o���l�<,��X.\P����s01)	����w/�lƱ	K.M\�������i�L�fe5���1��]ʾs��k��
�����.?՞�n}�"h�����_�I�?T�]�А�l�_0�V7/;��P}T�r~kc����=ׯ_�qs+���w^d�@WkQ0�G0�Ccm�k��-Y��M(V�:�5���`��W9��4��'�ni��z��])��N{#���7:�������f6�ϩe��cf]�U����y��#ͅ�����,T�^;�&-)IwP�����kӃ5���"��g�^TY<v^��&�`󰖛�Zz7�5�F�y���v�@�3]XPO�_�� �8���s�_�m�JP]?�:��Q��m���|�g8�({�]����qG�I�\�-begFh/o�R��lV��{߱��_��w�� ��t�<'�015�����C���c���1����Iw]��7~{�L<�ϠKԢ��j̙��&�K}�ұ���cTt�?~�^�)}�'���^Q�r�� Ƌ��W���I�<&����l9��'��4��98J,kL��Cid��}�mIs�>������z��UW�X�[��[�\��0 3�˰�T
��4p��4!~�{���ӽd�h��T�=������宗�0>�,wǮ�VM-�"ϯZ��m�Ai."����\o���a���̸������遪���^^�~���}��BsWd��\�UI�
���W���NRh�^M��I(�E�4��m���[�б,������YJRj����&׼����g��&�0_wIX��ֶpط���_�~��J������~c���B|tH�,8�ͪ̕`�K���!{Ҥ)u2\�}T���^^���͆�S�^�7�+��<��v	d�Z�kd���d\L������b�;��8��:��Z��.O�p���u%����:���8���G��嶜�����9|BBZ:.S�n���g�|}\JʸoE�9���B0𷚕���������\��:WJS��oF_�__Q�<ޑ'����w�F�r� ��'>/��i^�Dp�-C_YW�CCCCPu@�ˤ��� �m	��k�����L63��h�9SUU�j-��3Q
5s#}y��������˵?~�E�ZZv����h��%{�P��ZOɑK�]��*��1�Wݴꨕ5,a5K�bfb���_9T�F��v��ٌ?������ O[�Y�3�~��%�k99�UðW�� ͪ��)���n���d.�cP���;w�(߼ip/��Qx����Ø��,*�X����"#-\��V��f��5�r���K� �P��C����{�/�hZc#��sr��ZGld����C,hlm=o���������ч���2�-����̖�{��,�O���g����q����))+�4~j���}>#�;z옾��:0{iJJJ����+�X.Tȴ����^;<# @�4<���^Wx8��e.~~��勘Qw;�z[5==}����ϥ�]111����A!!T���){����Ћ�k+ν_7�K�Z���=�t�@�Ǖ�Y��gt�������q�'N���I�X\�.o���Cv�M�|�;��<666���T������}8 \MT�i9v㚆�j� �p>�`\Ѥ��tMu� *�j�/����,���O�m3��_�~Uz��D�QY�}�����#M�?���*$2��#����#:`���((��JE �Q����/6.NZS3�nɸ���^]Ʊ8��H�����sJ�B~����~.g�S������ם{~Lt�:vu䘅���T2��|��?z�(�[��I���c?��S;��g&�eT�Z�hWx�K��G�z�4`'���(��e[$VHXk��W�<e�qzɅ�Hk��
9��k�A)�%:���J�틋��c��؞���U�n6w�<��Me��~�*ЀC������8����Rw�DK�v�n4C�8�6��I��6�U�:k����0���F�D5


�7o�w�M9z�سg��n~� '�X ��wO]�l+�Os��}�F�͈?��ys������2vsc�c����h���Q.���^+�V�*ڻY-˟�L+��*>O����Y�s�xu�k�:��,Tڎ������k�o�yYa�X�G�����J��[T��v��Ԫ��aU�#b���ľ��%����sk��� ��j��M����r6Ϣ#����-"��������3������d�Ot������ ��B�!�j�jPX�S�(��fL=F��3�7C��$kp���kihm}#׼�C�Stlj���N��R�JikGP_v�aK��AduF8� �����1�6vv��Ƣ��T�C��~����/{qoߞ�3��%%��(�T392�F�P�`^GJ�K��.y���(+=	�����<+�`+[�Z�V�ɬ%�ٳ���Dv���#\)�^����\Ct}wZ+:g2��S�� `_�����|M�ݻ���|���BL�'������n���_'U��Pǩ���<>pEi�K��\�w;99 kI�����(���������O����%HQ�>{��m�W������?����G	��F�."R9�3F�	j������@���D�&�t5��Oް���3�����x����'����$|i�YE����#����@��q;fV֛�$���O��Z�����5��\2kMJ��Kd/�A�k�ƒ�-T�����Xnv6"\6����=q��ƦPAK_��˵�)��0u�k��I�4��K��Uƃ� �׿���Y(+�JI��ʮ�&_`�C�����<��~��5o{�#z���m���W������z//���긋�^��&!%�`1��gy4+�~U4�j�4���� u���H�`��V�Ee�]�U>���}�)
��PơP&�oci%�O�<3d\]]���]kL��'p���zS����3� !��=}���$`;8���nl�zmuYucM	:��L��)X�=��n���}��S����L5�.�<||,5d� b����6����Y�P��Nti��;!;97&%��.�ɢ��=�
 v0��	^!�̕�::��̖����ۯ|�v�<�vG���s��k�����y��j

	��@:͔�;:�F_�6�-��y�QW�mImz(�
�Q��}Jb��}�Я�N�za5��{5ڥ��c��n�}�̈́��`�WƎG��,���#�in��#4��������R�V0��e2�K��3��ebf��OCNnWs}���aee/��\*2��آ"m���V�r��M�u
��6N�̶̨����&~��Rbbbj�(��	T�{B��'��>��2�N�XER��c��S��Ԕ�Πՙ5rrr��Q�γ7�F1;�~J�MJ���
T�(���Ww w�i㛐J��8	��Sv��<zcfa�pf?A퉍��iT�hZ=-VWZ�ȼ-�����Fh�y�;=J.<xP.��hd�e�C��<����v�st�^��'TR���#;;,�pH��41���qT~Z�L�]5�1ޒe�#�8]uu��2W_���Q�0w�(y�W�}��>7z��DY��:��@`L*��:i+X"��--j*���}
ge�x/]���>�����H#��C�y�����'v�[h�R�&<����+�r�̫����?w�f��0�+��I�c�a�A��bccQ���l0k�
�;� 9�fG��h�U�Bvɵ��ˣ�t�N٨b-�F>HJ'�Ϋ���X48/�\�����$$$�uVn*:N#q�W�� �Cg�x$Nu���jv�}��G��,\궶9�dس�Y�X���Q��I��a����|�#�(�;\5 �i h�n�'d���F���T	M�E7 ʹ����C���nc���R�] ����N���K{�Ẍ�e>���7��Vnj:(���������\�\k�. �ƙ��俣='7zt�j�=��|h%$$P/+]�1OҪ�z������O��m�mЊ/���'��(ϧ_ �t>ҡ/ߌ0]0f"6�����
���8�ۀ�/��R���p_+D�Д���z�P�9 �E`��9�`��Weu����_�~��NH;.�$��P��ǻ���������³�ؕ1��_4���AtX�5٣�}��U���K_������dڻ�2p5�"��*�����#�������ޞVIPP��`XWWw�瞱�YK�R��������ႮT�߹�cAu�ȹ�-��3� 䢤�4�#,'*r8�ͨ��Y���0�eH�)�,��IC��Tpֶ66����9
�}�����?��N�����*)0�L�ˋ����Dd�75Q�.jĚn�Z�	�6��n�"�jdQ�Ռ*�����m�F[d���W�����EP���t�Rs��"�×�Øwb�@�р���^��n �{�������?���Ӏ�J*��4e�d�Oꀿx�6�D�[�,N��m\��$y:�������\��o#�G40`�4���V�El^�:j�'P��Dʣ�O�7�E����X{tt���T'�Bd �*Wq=���?�P_��CGtM�����j���ղ����D�$����d�R�l�v9�Nȓ��2�m�:�z8�S����7d �QVwQ�.'����A�L�
��N5-�p@d�A�5@A� �˅�]|�M+:˂�93h�o޼Y��L䣍1�������~�(�'��j�9�������ݥ�x�E2���Aջԛ����╀,�/�"��vxf� �tt�����Ɉ�
�ٍ�*�#����ظ�+�vzD�]S�MI��;~%��h�d�(Dט�2ס�P�с�w9}
�r�HS���r���$��'>�����0x���U)�����+7P�)؂@�q:������;,�	b��҆zɫ�R��)��Ǜ	QcD���˖7�����Uâ(�/''���2ps7)��ADJLJ2���`�ߝ�����b��.,8�
٧"���Y�O,,�`��� §�{��(���ruJ�~N
�����7���؀~��B
	m����
�~�K hp=�F�;�M�Gt�*���������cdD9`�/^H��D6��;�������Ld³�����;�!캔M-h#��&����R����p����=�U�]|����3(A�~Htn.���|2:$@!B�q�>*`i�aXbA�ڂ��gJ�v�=�}c�/��'o�H�m�� ��vR_rz/�*B�]��c����Ҕ�R[[�ތ���:phȨ=�*
� 'O��{}.��7G�4�H�ZZ���p�|���/_&�T�r#
X�Kߜ�jH�������li^����b\�܆����딢n��礗ѯ�*��?z���~G�ӓ�ϊ=788|�:-1QyԜ�u1�����2aM�E��O==�ƿ�t�+$�4Q�t�C[�*P������*�R�͌�=�lUUU2�i]-Eyy!3l_�fg+���6z5�s���ϟ{�,#��h�o�)CV"Z
��>1��3}��l�9F�Wv(�{s/���K�8�<:�ݑ����n����~g���.�Q��AC M(�_~�4x�عʯ/����F�
ߠ������� F®�K���,���f��
�Nͻ�|�~�ɍԏV�TƗ6,<%Z��uq2��虘����e�����������aQ�-3��h�/ou�~k����U�
���Ӈ؟x{�1��z�/����sѯ~ 7�GԀ��]�`���<��� "��l���*��Ap���?�@@ښ�j�MAW#�	���k+�(�x��F�s��Ͽr
u؅�[_uu-b�W������Z٢hWvũS�]��7wEܻ
f���ăv���&� �f5tBQm�3β��9o�K/�����\�b�qth���R{��)d:͙6�M9\F�D�e៼;��#g222��<yf�2}HZ?5�b���9�"� B+�4�1����:���<id���ړT\y���%%�^	��r�;��n��⽸�DVo��� �eHY�اϞuM]c!SYt�����LZ�hogՠ�O�!;'GZK��m�UPPB��3�#�	��+Q�+0�wOJ�ݽ'�%p~:�IKKl(zWʾ}���\���E�����!0$i9��撒�ռ�qu]2	���%;]�[2Y��f�l'g�4g�����M]�ȩ�@S�dkKqC�[]S�G�ܙ3WѾEʛu���+S_�AV�A�Sb_Q�$� �eYg��X��h�Ց�9�#/6�)^K��q99�0jՐ�H���mf=T�p<A!BY����!�K��O섧��,MuTU�>m���(E����ߨ��-HZ��r���Γ}����6�O���?��ŬC�B!�D"A��0���=�ɍ<���G�Ӕ	�|`eq&~p�Qk�8-|#�@s��u��K��{�cm.�|��&���ƣ �!8��paJ�N��gf]��5���#_��5�j��b�;�u��Ϧ�ڃ�y�䉠���<fTf��nl=,O�������>@��?�F��5Ͼ���Q�6��/��|��#;91�%��Wz� ����{�"�T���6?�y�1���D.6⍯�����+̗lh��G&�
���g�?�9t-5��1--�L�
�M�� t�T��gi���e���`�߽O�y��VY����yӥ0�L�?u����XZ��������k;zSZ^��x�x��s�@r�᫬;��3MOSS�
�ֻ���y��7$9t�%6q�|���u� 8A����l����j�&�θ��n�T�DP���xCW7*����GA�>D�����u?��h��s-:�4�7�~dr��X��ݻ<4��o�+���H����&��� �Zh��� �����~����_Q���Ky������V��+W�E�F���W�'��)�{�|�u���2��.d>1�IP*|�s��f/^cc�\]W�I����y�	�e�"����BK2��yw9����`6�KY�g7��ۜs�6EB2��
K"��$-Fy���t�˓%=��+f��"�����&|E������[�5��
'F΂��ܴ"�����P�T�H;M�ay�C�JD�&��2z�����~�7��S�A}��+z���܊ѡ!+b���g�N����W8�n�+�|o���+`{�ۺI��N�@��q"h�����qB��|G���f�g9-��@��d��"��Zl��e���a"���<#>��m#D`������x��c0� �^щ�վ=pN�hx]|���L�z-'=^*��9�D�6��5��#�w�R�+�R��\���$4
�R6�
�v��I�KN<������{�����
rپ�'�#��G��f�A��cK"�k��&�6N"�Q?��mλ�x�B|~��R�`Y(d���`�~�Pp�i��_��ZH�����G�<����]iD�j?�ٳ(��}}wz�^���%^��GKA�I�q��J�ߧ��ʪ������	l$�&o�D�{큼�m˃�%���zԴ�Us����'�Cr�%�:���J]I�G�J悋Hs��k�w�}����i���v�����XKJ *z���x�|��v=�>-#��v����x�q׼3��
XSS앟*D�D^����}$�t��y����_����.<�x�����n�u�F�S[6��yo�ޕeܲ:�A$Fla,�2i?ޓ_�#-���Z2&<�n'�3V"_�+\�ڊ7\)-�gQkS&�|���'��PU)��[���<f�8����+g�S0Ba��|S6������5��$�A�b�O	���w��<u������t��u�fD}]o�덚�"q��{�w��d�$�IB/	��v[�L����z�!J���/짹����؏�k���n�=�s^nƪ��eE=��R�7="��ĥ�X�\��*���]�Չ{\B<�w+�Hd�LNN���g���ّ���z7^����_�X�}���2���P����7�@PŠB�a�u7�K�u��N�p?]�^b�(_O�����8͔ܯ�'�۳	q
	6ŭc�2ý�α�x�P߯O*%%t�#]����������5��<��]�p�]���Ox��;���/���SӖ��ق�ۺ_���#sN�^*��G=
<6PE����8�o!�g�[�Z�DA��Q�����9�r	M��^w��Trm��.t.�ki��P�\��j��Z�jKީrr|CZ�j7�ͽZGoh>���0I�F�f�)>O3���A��.�x�-;-���JŒ���x�����1��[^��޺�j��5��\��	��NTX��z%K�Y�ua������X1|�u�B�ֶ�<����Q@�j	��nYס��{{v�x�����ۮ�¬O�\W:.�H���-��
��Kwh_h��E)jBK�0{j���vj|�̏i77�	�oa蹳�*���^-��YId� �:��c�|��D������"�a��-��֎��&�%���j���Q�'=*�`��!�Ԯ%��$Ba;&M����]t��x{z�4h�@�o�Z'5W2ț�~`�Y���Ч�ֱĄ��!?���\ ��P8?�����W���	�B������5��*�n%Q��_8����PH�%В 9<);=₷'��.��m�MС�wt�B�/h����΍��_�W��0VOW*v}'��mW���x"E�Eş�|�t;h��:iV�s������OW͝�> �a��ӣ(�36�Ÿc2]��]��.�9e3���8+���Ლ��~��$Ey����]++��o��-�CP�n��A�Y2��&�t\��Q�l��2��.�1����v�C2�|����D\�GO���k��j�W��|x|uk���]�.�'� �����"�tZ���.�.��Y� ~�
��xv��W[|�x�H�c��pd�~��o_�P�S��U�<�>���C�i�4L��咨ӫ��������far}m�_����X�5!.�d���\������@�Sg�5������7�����̲z�3��s���P�����hz<�O�,|s�>&BwX��U{,����X1��_�EfB1����2EP��v�s����\$A���s88�eɷsX\�1�������k]���y{�:}e�9OF��յ�RH�*�S�/d|���X�LD��IS�=�S>vȳ��v��d��yfd�0��[����S���,y')i��µwh+S�
��2�$v��Wv��\�l��]�<��u�)��o{�ҏϷɨ�q{c�F\��Gl���sN���Yk0Sw�	ٳ������T��my�L�,������_C��,�ȩCw���C��r���>bC	AΩHǦ�����P�o�Zʚz���Q=ى��~�����������"f��+ ����p�i����tI�Z�u>����Мs��N����*s��Z�6���ZB{�C����Cf��u���$�('v�����'5��~O��'M��\r�)xE������k�֦x���sIO}�Z'�(��>�8s��L�;YNڷ����|��)@��ǮǼa���{ܮ�qG��n�Q;�Cީ8�П�r�_��_��.-���2	�-�Qt[�l�ۿm���ދ�1쭴E]u�����
O�L�yڶ����P��Į@�w���N�8P�9���zOxk߉�t�_����FU�n#uXyy���1�*{��b�6�{M�x�ެ>��1�����
�_�q�	�s*�B�&cz�;q�I��'����Ho,��PX��s�����t�Zct�ڂ/�Y�;))�UX�(%&V����a�~�e���B�ֵL����=Nz5����JX�2:<�R�V����hZV�ey>���K��n{�t�/�ZYM�u�6��܎����p|� Z��c3ZY���O_|�>�c��\�p�Q��a���*��k�}64�/^�}»G����C�4�nw�����>��Mkf��1���la,�1O� 9��g��U��F�V����=������x�*�gnZe�:,ƙu�6�$�}��I`�촯��]K̊��1jI��y��J��O0��1�3c`Z�v�;�Y"ߺ�3�Uf�_�e4R��8O1D�툹��NE��N-Y��l^	��˄���{��p1���߿������~�a�,,)�:pӠC�o0�Q_���\�3�|9%c��P���9�w�B��H��u4';��qvv���	�"M�qxt����4`�c��"�����r�#�z��; P�g`#c���w�4�k��ou�G�	 l+�⣑�������eE�u�Z1ۗxbyy�5�� 櫇����~m���?�0�iV�DwD���#q���#�J� 6����S�*J������7�'ژ��wk�\9�Ƃ�9�X�X�������<�H��9��&����잝|tb���Z{t���2޺,]~�3ֽk�$��d@H3E�9�d��u�,!�ŋvs5�mW�/"��N�*��3^57��/{΍�	��p֭���ʊ�N�6µ��Y�3W�fn�N�]�k�.!�$��'ꌸ��c d3ͥ��h�|5o`��	�H �]����T�C+;JT���fwp����@���Nh)��!߽h��9)qD���m����~RX�=�8q	����ó�W���\�7i��W��mrN�hSS��c
^Ẁj-���)�����+y�z8wmhž���V9���W-vZ]x\��|a ��L�Dgҙ�L�Np���̴��{}�@�`���X�/��2���,���r���~µ�umCXe�H�����Na�8��}H��\v�t#�<0�Z��д�Q�ڞ��zM6uc��	qu��>��[�"�U%!�9Ղ]�FlLVQۚ���b�E+��*�L��mm�I��Ps�(}�鴚��v�t��~�|�o��Ǡ�W���{���	��}̐�R"�����փ+M�X>���j����^6Rއs_�%�f�G-}��Zm�J�G
����KZr�1!���n��l�����������ǳc�27�eF��da��~���]�H�(�1iW��k}�0t��zkPjߒ���>K:"�t�*KJ�A�;���N�bWWW �����>�͍%���qo�[z�q�����7�٢w:��D�`�2=9}h�@Ȗ�ni��L�۶��ox9���<rD���z�φ��<�X��_�8���f������Z]vb�0y��ۼDӚxs�iɲU�}�	�d*�s��Ic*��/m��Qʝ�'��x����8kV�Qʦ����3O��`^�v:?���*>,D6�s�?uN�	��3�G�������ϻ8��)��&��[oӳTw�q��2��r��	�I�^S�s����K ��!�j�Jxdk��9��\b����15h]e���N���@�J�]����ͨ}Q��/]��w�����e#�3bfS�ϊ�bs�t+��x����5�>���P�g�q`ZŢH�mң^Qa�S
6�u*J��^o6��hً�]�Ou⃛j�0a��Q��'�B\B8�d~۞��v�1cs)elAnt���~O�D�p�����Aj��2��7�x���r]���k��%�������5WD|7��������L<�9�u�C���,��?���|� e��P�:�6�7�
���"�ܻgvd\/KS��</���/1k��#�h�Ԅ��u��_�zy�NX�˰l�,WG�@4X]]�)�n�0nPҰu��������};�lnط� �@46����KN�WK�����n|Z���Z��4��ey�k�����%�|�6B�W(�z��I�s��~�6�N��p�qSc��m��+����U,�z�,EJ.�ZD�Xj�=�S O����o�v H�Gu=��^�O�Hۣ�}+2׋R����~���n���T4a��N~`p�����@�z��D}=����P���9.��<Y$�"�>r ����*	
)jB-�[+��,g,�6���`P�8�?9�9哝T>ߕՋ�r~kr`Ҳ����I;V�*��3\�����E2�6��������T]ӥ�ݮA�c����:Rv>��ZVH�t�F�Dn����e�H���Mh�..�p�rx7��N/]�0�|a��@�������������:��U	/�90Z֊|`J�k[+q��r�G�4�Ӱ���	xϻ����znY�hR�w�P[��O'�d�f�ԶeX����=��~��9�g����B��9���m
���#�����e�7��s��7昼䱼��6Msp�qN�L������Y\ ��#p%��Q��%_p>V��O�+�@��?p��'u�m<�96ȪrT��,�_��ʬrV{m�Ј`�B�NZ�Ÿ�����I{��KB��2�J�u@&�>hR
q����	q����8ֈ�1���m�����_��Y�$Ľ�9CvLy'ѓ���rys�[�s��ϗ�F��1���s��k��m�+P%jcH�������ez�%��W��^�(���'G�g�Vߑ�ƃ�9_g�T��l]��L�|ڈZG-\P:�R�9�)��[A������L��z���&o����F2��Pp����[1�W��Q�4�)����_�*2$��I^&�f���Ϡ0:�b��q����h.��ةnS��w_s��z��e�C'X�b,.��u�%z+J�Z�E$\�'%#����ms�楡A���j��?,~�~0+%.����d6��Jj	qv6��9K�nr	Ml���}��乬���xI�&ٽ�e:J��m"~S��������Vrv�����R�:�����y�H�Q�(��?�?
��z���pWY�(��I���5&�Js�A����/���V|~_[�8J��9���n���Jg���a���[>�3��䢷�.BP
�D�9���Ɔ!���.��n�� ��f;�p�R�h��<���[�Rd,�qTJE����Iu�>u�nM[�H%nz͞��"L�E�ؠ,��'T.��C+JՊ-�
������\�`���Oh���"���łh⏲K���	qn�9"��m5���z7�;3�mV��2{=��u"cc{�6���[���]��Hq�'��� �����[��6 ĊI��{zz��}@TQ-Ip�N���xqO�	r��P�tt���k�zƕ�Z�eS-=.@LT��S���=�UT����j6�L^�"����Z�+����.�>��-v�;	��𓩥���s�Iq9��d���߸�sp�nç�����M�"�c?.񆙤F�oN����]U�ܲ޶�~';J�SX�R�8��YO$���1F����uX���s3z�34+��L�=��	���1�=�E=�ea끏�X���?Sѹcç�q�lE^��s�)K�2�8ۂ�!���C�ݒ�e�1��zi�#�Ld*:e�E'$��p��@t��J����[��8e@>�a����z�Sg��^��\P��u����x���\����T��+�%�Ȝ׶L���G���Ԥ����Qda�����iI��T�������^�k�͉����7ƴ���T�����-��w]��n`�o�:9=t����1qʁP%))�ֱo`���9���ͦ��r]��u�����|�_c���,�^��	�I��Ʉgo4��h���󹕧�W|_ ��֎2ɝ�@C��&����'&�OLX�����TԖ�t�2��!K�o��U�͔j#	ӱ�tI	�f�0�Z�k3ڦt8��\ה����ncyn,k}k_>�˂SR:~��/@$���\�!�K
���Ӣ�~��}l�%K�oy���W�W�=$xd�l�E�ذ֋~)���9�B��0��h�g:�?`�q.I�����予�{Ii
x^@Q2B?l,��3�b�I�g�����XR& 8|���]�͋U�O;i]��������\/_<6�61��^�f�2����,۫�'����s�N���U:����el��Kk��?O�w�����AS����S�����O+ ������籬�Y�#�}K�0��,P����OO���+E�3Ru�{��O�s�ñJ6���퇦�'���S�Ñ��Pl���G������I�Hu�⺦�K�kL�.��Ңm�������|��p�í{���Fj���H����')>��%I��[eE��<�/ �; �///�O�C��\���s�\-�.��Cr�1�g@�/�|p�i=J�X�Q�����v+���s���z	A����o%�CE�����0�6�����W�P��J߲�>Z���W�B�1i	(Σ$�D����Xݾ"�w�n�S�&"х��j�be�CfB\-�GeE��Oc��\�K�g�^ק�6��J���R�L��l�0y������s�6�;e�Z��m��F��.x��"���F�ǳa��ʹ�l|�*��\;�[� 2�i��d� Q��iSy����I�ʲm ��v<gtpb��Z�h_Ѥ�U�E�4U+g0��V�}�*+z�z�@�HĤ�q�L�d���W7��fe��+.c����	q���&�{�ܗ�ܩ$�n��|Huh�f�0�p��?���	[�,�PF��n���+j�Wj{ `�d���:�R
�;��7�ӻ��}B^?M�t__�Zj-��4cҿ��j2�yi����(M��b/F,��c�M@�����Y���uN�7?+n�F _����O�7+�c��r�SB%3BSݸb> �����a�)�=�M�o~?9�y'�|��\��ʐ՚Q�뤷e��-C�#g#�h��>��r�����èl1��~�I�PӕŨu���J�(��/�Ifh�>�ϒAE@aY#���6��f����32�Q�?��GR�ן�a�]0���6+��3Q8��:ߑ�[������ ��MJ�ŉ��$S�d��wV<<�>�p.�����ML�L���}����L$��a�a�}�}ɿ���1/����zzD[\�U��o���儀�4��"�^&�X޿�AB�� ��b����w����|u~e��ly��B	�c����M����;�N��:Q>��{یл��_��i� ���?�c�^li{�7�c�hr�&/����^s�7���������rC��W�M���3
i�4X��1-�N�� ��Ov�s�w��<X���( �,gZ1"ܾ0��d�YV�U=T��(_��z����ۆ��S��I���
 	�Yu�j�]���q�u�&��A��V���x�����;�9������țo�F��;3ހ���� T������T���J.F�88Qz�	�Q�hMT~a��N+�5���oee��4W͗s�����;J[<�_A#=�⽴=HA�&#I7;Ԛ�di�8=�n���s%�}�V����q���ێsN�G���N
�I
Z�G���3�*��Fi��Ɛb��o�'&���"y1�z�q����z���\�Ҽ��W�#��j�s�St�S�3G�����;�h ��a<�+�1�A�,���޺+}�&ʈu����R뮎��8����P�R�LW��.�ř��H-��5�\�N��]t��_�����:��=2�<�Ҡf���:&��7�Kq�^y��F9י�CE�4���m����/#��|��HD��8g��hF���$iӌn�^�i�.[�¾io�jQ6��pڹ��U\O��6/M�1��pu��� (������5�����{o���;mN{"d��Y�C�,�Ȓ=D(d�`,�S��첕5I��e,�2�Hv����`���7e��{�}�|���u����u_��z��{�,�cg��S'�fg�f�I�����30�WP�IOx�ǃ���k��z@G��"z��?7�L�-�B#�0*&k�DJ��t���v�|����=���V-գ�l=R'�h����7�����á[+��ƕ#!�÷�=��k��壺�p%o W�]���IN���D�N��n�{�lMBA���:�^u�������g�Z{���X�����:c���,� ����\y�I	���χ���U9�� $ �Bx�U���`{�t�#z�cYy��G���Je�[�n��g��,��*�9RU�2�i�Њ��[���C5k��#�fLкn��;Mߍj�/0��pn:t���6�l:��yKq~MU��F9���u���&mN%��fn����6U���7�Cseu��a4}��̀ùa��������<Ӝ�0����f!�svMǘ��c+��d���-.�I�eyќ ��ˢ�pk�aO�˽8BN*#x���[����>3]v
����<N���� (��������`��d��G�(�xi��i^ʀ�0�@�<���r;�+.q��L�ҐT�W��}�8�T:�W�ѫxѺ�И�S���Mo�aR��n&4��*�Lw��Ob���;�I��z�왹W��3�ND�2�,í�=0���	���9ߺ*�W�6��a(�c�
b�}��~��Gn���;b�}���A;����� v��������:v���.������1���Ď/�
�+{�4�$6J�Yl��ОI�p�"p���Ft��t�3|�2́�7b�ȸ���yod<u��&����q!�V9�59sj(l<m�e�tF�l��lI�5�m�Zo�fߣAl�WL��)حz��ϧ�>��'�(L*�}L�����i�q�2@���������?"������P؛8�\��� �k ���*_������q�Us���ה����o@�&�Y�w�v�򤡉;���K��*5���=bV�2S��<j��=A@u�}J��B5��HGUQb��ytZ����W�d�P,P�Y!��օ�T� �� #�5}�\m�m$��:f63(sJ��o����D:]�����5(w��u[�q��^H�٘p��vW��s�����
� �t�ɣ��c�������պ�W��Fj���؞ݏD�A�v�:l=G|���c���� ;��b�c]��0t��E�Ƒ�~�\��������E�x��w�=Ip����?���'���v�a�qaa�DS�l��k7�=���sȉzH��C�g��8�d4v܇l��(_;�J�5/4c�QJ��se2\AK��������h=*<K]�&�R�sGд���!�h�(�x��tZ'��g�����%q|�?��9h5���v�6�e5ol��b����,���y���W��S�5�nf��˥G7�:�u�y"���g��������zO�9�o���y$��/����۵J�M��D��wI'�>e�/��4�x�_��c�{h�b?G՞v_o#���p�-��+5�?e+���\X�Dy-'	�$����+��#����̟s�=��eE�|QQ s?��UՐE�P��;:�lu�<!wWS^�����m�o�G~�*���B����0C��17�o���<g�� �إf���qAx�\�?�g�0x�O�Z3��c���~h��wM��.WK����!���ھ����.�<�t�#��d���ܽ�{�}�)��z����KG�д�l6*��B�d�'J�)j���k4/��br��1V�;ހ�c6Fb,��f�P|��}�Z���]�6J�ֻ^0� ����J�Ll|�5������H3Q��\��1�>s�Hhw$
Q���6�uw�
�H5����.�9��A��|�Bp%y��:��"�#8��=+9��q#��"��K�"�MO����h̛t��Dl��l�Z�y�H����9��ͅ���ê�B�]3��c��~��&@� �C��i�L(��b���F�I٩gC�_
�Nq9X͹��_�*O�Mn�zI�17,^�!��B]S�lk���7\�������cG+y"�L��$���y�	JcT�|b�C��M���+̘3�cr��T�qr2�0�BPPP�j���mFp�Ln�m�R��	�+��ݜO��ZYM��(�̔�h�!}��g�^�{O|ѻ�V�$/C�e�l�I��Pt���S����?�8[F��H��ϋR_�����[�6�<4Z�`|X�h�u�AX�	Uˠ����,�4d���Ox����Za?��uB��x�˪�����ǩ�I�.R	�:��<(���/%1�!���������+ۧOW1�O\��^��H2o�2�N֩H��EEE@!�O�>%FN!��U�����i���b�-��Uth����b�{C�[��diDY�J�;/���ӑn������q�m��/Ck�&zФ��\)����u��#���[M��aI2N���tt[��[�#&��=8�TȌ��!��X'�`cr��B�Apvv6�1?��ݶ秀�lk̭hWF�]�;0]7�5d�iE�uc�W�xF�� �s��m�m�\4�Δ��I���H3��K?�
�����>$� み>UU��E��\��0�w�އ��y����϶�h�U�Q�Y�҃����=�w�NJ�����$#e���=ȗ�Ru��VHQ����k�q2di��'��ɸ��.� �LdW�6~,��N(�e	����;�>+K�"��}o)�E�.�l�����d>͖�b����������A�+q8Thp���<@Ë��Eu�
���z������/{�Nl-���E���P͝"7�*M�gr+*=G�9�uf\'�3DM�]�i�_K�S,�ty=u�ô5�S���_d��>���y��8�����ētt
�e�!C��M��#��x��js�7M�
g��6�d�'��D�T�3а�N!['� ;ʣ�рL+t��/8!!�9x�O��'=����)�q�0I���R�H��~М�g�$7ֈz&&������π��(a��$}YYY�<I��2]̙'h�y7TK`V��=@&����P� ��gM�Z�	tM��j�����%�°�k�:@ށ�1]3
��զ�z0�~ ���pŘk��ݗ�������_���I�8 r�r&�[2\������װ���	�=0�;Sd��ה�X4,Y�HsE�ϊ��sn�	�������Сk����k.�� ��~�{Qs����
���m�}�Q
.,��A#X���i�.���>ޢ�[�0���ٛ���g��?���<}�6l½ݺ�p^�e�6������X�5�w9Q��B�B�~p�΅(�B�9�d��L�௜�c+r[?��nC�����r\_! �M�/���1l�=����j���G`���Q
��
�6�:�l;�r�>W��'H,�XZP\O��Y������o���g�g>������b-��ي7�]~���E��/�>qI�%��W�X�]��0����#8@O^mu����[�[[�.�U��X�ِ�\^;��?�E�r�����Dܐ�΂L�LRg�(Vy�G�<����n�Ti���X+�e9%�˚�X��:f
W��l��aw���UG�,�ʥ/r�]v?R�4I>�f����8)P�m#tEO��fWK]�M_f��U`�{��pw 0��$R�b� .�d]7)0��"��Ͼ9����6��R�o7ͷ{��d�ښ��p庑��p46�h�����n�����1�>�߉+u>�%n��)U�|Zǟ<� (p����\�̉���KL�I+�r��j"��1�j��>z�P9:66��Y��"y�.2���O0�x/g�>��{�7[o��aTQQ����j�\�U���sk���Xp�֓+ ��_��7 ��E� .S��[	Wpl�h�`�0�Z4�.�d�;rͱ@'�%R����6�Z���@B_�]e����`h�zWr�~4��?�j�}�2�r��m�c�^��Ջ���D����=��Yp @y_Y�S������2��|e�g� H1���S��tЗ��v��ˮ�;t�d�P�!ϋ��M&�`���@Gg+a"ۓ�s~�}}}�Y�9 _o��DJܲ��g�z=k���+���N Dp�)H===�dJn�^U�N��$<�,O�8TUq�W.`kdy�# x����h�KrON='��<��^zt�?�D� �ĕ̫I͇��HY�Q�52�ѪBXOc~���TZ50\	{|Я���U�H���߂g���*NnJTǀ#^�!O��P�����,4�:�[ȧ����ewPϼz���1C�N�dHژ�Q�TF��'�ޡub�����i�����i��7��V;0l�f�>�WdQbw�tZ�>�s��D,S4~��QFZ^ 3����v�KՔ�=��%�L>cY��J4c����� ��|w��Hޘ$�sO�ѹ'*�i�[� �א�'x�1�Ve�ܤ%�P�h��ї�U��k���Dx0V�g�<�t-�u��� R�L܉�G��]ɕt&�GwgjT{�����QI!��IP��bƞ�:她�
�����k]�9�R�0<��ev"��gW�bWTn�,�s���G�#��q��ť���Y��55Ғ�����*�Z�f�
!s�X���	_q������'5g~ρ����r�8� ��y=q�@�#�'E� |:����M��[E��������\�{����������j1���pWh��X/�bo�uk�;݀�G���dc�CxLzn ~�R�,�F3�Z ��@B�z�!����疗8�L��f%qA�(�����NY,��)�k����H�}Y��#���ޒ�S�+}�]�N)��/�H2�K�(�6aͭ���]e>�u�ީ��}d	�B�a��R��y@.������1݃����<�6�L4	VR<��C1����uL5-�n�G6��r
R�����5���*v�b��?	���X�%4���yuJ�~�����?tt@�!�����]3W��ψB=��}r��Q�P��M�������5�{� �j!�d��2�RN�
⨩TU��?�<�h�V����2-��9`z(�Q(�p�>�l�u��m��T�W��/����L��
r�����qqq��@�ĸ�A���Alv��?.S�1k�ʃ�h��în����{��j:�Ӎb�&�Z�`ɜ&��BRŐ���[^ΆB�rKJN�thA�Si��Y�JI�"�k��t����QN;	���#�نj.���{���V��y��BFJ�Oʲޟ���z��!vŀ��d}{8Mz�pt,��'r%�x�X3�}z"e%����ܢ"F�Ǒ�`�kx�P��TZ�
��J����'6�(JQn�Z��_dp���ͪ��Js����sۗ�)���NKK��? E�N�{{'�v�<X6�u�B�I4 ��=zt����fVV<�e��`5�p�<����OXخ�{�`�L����X0��q������ɓb#��󛼋�T��M� ���G�#Wh�o���G)�o�T̿�~|��Cvv]}�" ��{Er�ͩ& ��M4�A~���NEje����!Y��z��Nq��m�6gs2�1Y��2�5�0<l��V����th�K�e'+׋9C]�o �{5r	|^��lY|)(�x�q�}���npddv���G7l�Y 1�Ɵ��$�gѾ���=�Dl�M�21�{�����5�4��P`@��KJ�}��T�X�AQG�K�rS@���UZ�A�N�RB{��/�1� *25�,�դ��g:��{{ �6z(Β��w���]�0�*�?q�n��!63BeX
5q���{(i������<k����;e�Çۯfgg� ���+��F��>F�9����XéW�W��B�>�l���͎D+��L���̫8�?Ըk�R�F��wvv���)���Ѯ�.e�����;22�A|��=p���99j�gs�,٘�8�z��ei��
1��(�C3�*�;�
�Ѹ*8�+�{mW�`����d�-,8���=�x2�TŘ뺰ܚ|���4�؅��wB�߻�`�Õ�v�H_7�W��I�&^�.KHh��y=�LL��Y�2^�R��2@��"c��s�mAJ�������(�l�o�C�E��G8H�"Yd��i��_��|K���j�d��
�b��;]a]�;vi:��D
��� �&d�>�S�����`<:������*++20(�*�Ak�����_ĠذS�	A����N/�Q�{m~ǭ�'�j���8����/��-�� �fr�*��M?�T�$tg�p⽸�_1E�ˉ�����BܦX�F��9���#�b�~�i��E8�k"-0��񸷡'��y��L��z��>#1-\�D������.�FZ��˸_T���6` ��"LL6� ������}�V�;��B�\��~�: �-���5�Jz��FzPiw���d��:���8a�QX:֓� [��]p���N�5O��p�z��F�u[6��d�n7�53kSBeY��6\\�zs7�d�=�,V�J�̊c�ā۳��Ml�$7P����T�<Ԛ�,?�U���W@�O���@����`�
'?^�V�V!��Fq����0L�$�f$z��5}�>��ı
b��g����~��Z�9T��c���^2����\��ؘ�r���
a$3C��re���0� ��fR"�72��d��`��Y
�?�����;�M��e!�@UHDU�9ٕD��R'��m��z��+\��;�BAG�v�����.R�>U��h1�H��P9/nbP���Q����˦���a�#xz���h��	�L��	x|iP�zP?m�⦞�͖��f�I*J����?O���j�9��Ob�;X}X�	�y,^�yWϿ��n(�n���99X�PD�G}-_ �믖ӧi��6�y͛g�a@V1�f(�)P+?[�K�ʥOkõ(�V�񰌹���	����b��z���"��x�8}�ϲ�M`��6pKD�`�qNF���A_{
�d<�K�/gz�.��� ��ʐ����yr�Av;=�1����e-�QiƢ��X5�4L��.+����Jt��U���׽hĔ@���׊1��#�:e!�Ӝ�H��8��՛���1lڻ}sAu#��B;\/�}�C��k�S��J-A��Nx�e~,��[��zL�z��0�Eݰ�<AxNW�7,������d��1��bN 01R^�a� V����Σ:R� A���
�;�G�S6	����8��üi�'z�G��/��Ќ��o�R�Je�!�;�� s�� w6#��cb��9âV��4�����)fL&B��2OP4�a2��~v��Zqc�<�i��$��B8ON{�;8_����333�:Z-1�O����_7"�3��i7˃�x���{��B__���!���d�O��جd��s��T�H3#�ܔ��K����aNG������z��7 ���i���H���o�-3?��x1���n��$!�
ӫ��,��g�v$�՛�󪄳��W���Gg�/Z	콧��������=!��{����<��,��ȴ���=�V��2Z~c+_i�*��XlP0ڽ�����㚓~�A���3�.gі��-<*>�v�k��>#]E�n_Іĵ �%Y�Aa� �h5�2���qA�0�V�m�׮�ax/���Ӽ��wr�~�]��,guP������G��"�s���ey���Pʢ�a�5��q�~5����M�ʳ�aJ�:q�y�\��	�sj��}s���8����TE��m1t˞�1RT�Jk��_th�27�pt��3Vf?"���VjTb��;�=WW����U�ע6��>��`��:Ҡ�7|A�u�� ��J�3ˁD��D߭/��bCL�/4�����<�SRx��B��m���[=��O)�O�&)��oWx�64�^��`�ts��)�m�u�4gN��R��IU¨�>ǳdW?2u}��� ���"..T9h�LƜ�@��I��!�[x�)�IS���{�v�mj�n�It�Q�-� �?V��q�)��}��TB��~9nu�$�9u� oG_(l4#�|�� �T���e:�q1��۞v^���f�������Ey׉�����Y}�$8C.K���X&V%�X��C��� P[�ܛ��}$��<e>�w�	��#/�jHe��'�� ��#�)�)2�6�#y)��C=���"���F��=1�7H���|���r�-�Uk�{����9j[�r���G��A�J���g	B����{ƈo�j(��RT�<��g��T������ UJ��*A�#�M�OxСy�/��\5C�%0������b=hmܾU!��P�Y�e83#1 �U�<3�FN����$[}�a�pZ�q ��CX_l�:� �0��C֒���,LW�R;yU|f�a�T)W1O�nN�&��.� j?B�r�b9}d�G`��k�s&d�{�W��	�<��C�'g�X��nD���F�s훟ٽ{C�=VI�VI^���˙��GyFJ&�k����g�,��:�5����d�o�$d��d5�Ŀ�s\�`XI4�/򺗧�0�����0P�����������ko�b��Zd��eW�o�.
���qA��N���>�����a��P:p�������Z�8�H���u����\Nr�� ��ۋO��<Ɣ1;;�.g�7n�����Ü����Բ�:Z���v:Gպ�����&&5�}Elr�2�]>�����G+՜�� 9x/J��)�h䱟 �y����>�	� K���.|>��r�\�E��r�>}Ɓ'XØcEޕ:���VV��Vр�i���¶ɐ�gZ�L0Ԝ������j,�~r�Cn-(<�������r�666�"XxC���p�)%U�% ��!ItX�u��Z1Z`��q�8%6���l��hӈ��>m?����_��ɀO�O���vj��1v-�d[��L+\+ܥ��1VG<�������'=�*�U�7�	�n�R%�^ �I�0��pu3����f1�^�PY�0�O�*"ȋw�D6Tǩ�l������j����M�Ζ?rOD�W��u�Wx_�1澿��:�y�+��==�\}��yY��'	���}?��p��r�Nd���W��9処M���u����G��W���ǝ�7���cD���Q���k�M�'�̎���ΓQ��4�ZY81�B����o��A��(W�=��B�I����`X,���;9?�n���X�<�7� ����]-X�q)�{)�4��Չ$Ι�u���o߮�o�V�Ux��IZNO�g��G��ߍA!��f������cU�v�[)�vT���mi�\�&����:v$���Dx��7Go�u`Eq8��K��G�^��>?j�U:�R���Y�71Ev���B�����N�͕L��s��%F���U=-3�.���r����frPv���G�Ծ��ur~1��K`y~@n
�Փ����-����y�/�(��qb�R��Zf�T�*�i&#B8�8�V��K��ᭋ�%tt�w]�#���kĂ�T�9�wS������s������ťa��m�����|�B������Q��%"K�+�i�ܦ��@sȒ8��ߩ��ZK� af?*�s캋</%�e���%ғ/�x�f��ѵ
�7P�D]�Y]��i~�3C-�����U:��$o��Ͽ�p����L���?״�W Z�f�f�IP����V�h�[�*�1M�*�/�;�v+=�s������- �[�#����;����9�9���E���Y:�Y޴j����E�]q:G�P
�UPa���L�vPm�wl�	w������XSS�ObfcS-�6�U}�+kY��)��Aa�)�����p1+�JAEjmC=�hH��������p#[G�\	�ܿ2<+�U�F(�qS1F�� p|�{~���Cs�?�U�X}��m!օ�lLN>PUUM�8 ��ݰ0b��w����AA����vl�o3a如�:�����Y��?5#�<���C}� �B��������t9���%��+h�>��'�z�*"�(������1 � ��`�����7�Р�)�|�iJ W����,�\T�j:Uhp�Ճk|�H���Ĉ?��j@_�O �m6J��Uu�/�v��w:Y��h�.�(ׇk�I����|�U�� ��M� �+��h��fܧ&J	�*U�j���ϥ���Tw�l�G*� �<� ����o��\���I�\��u��0B���c+#�a��|D:��#q�`��'���*��v�t!S'����>�1��D���h���sP٠4�
��oObm}wN���/Z�Ui��q���}������(��hĲ���SZ���/�:����^}����{��9�4z�	Y~������V�a���:ԦH�>9U�$�10�T� �ˋ�i��v��}�AY�q����sgϞ>;�t�߬�S��Ā��-0�o��&��^x`x��3@�e=u$sM���ʎ�zw�~ʚ�'��Y�3����7�H�.;A������0S��4���<����zxQK�+�����`� [�98פ���P9���#���o��������R��W���
��ԉE�Z�������+����%qn'R����Q�����m/k�XWt�w��zp=���;>��\_�|C�6tƈ�;�XDM��ng��u�i��i:�h��/�쿝�qr���ƞ�d���W�j|�A��2({�bص�����;�x��ʉy�NLd�x&= Xu�������3P9�x�����i �RR�ť���q�(��=������q��s�v�1A�K����M�f��)��I�8�}���q_�"����Ix�l�`�e�5>r9���*m��5�.?�G�b�{���K����r�,��-�{�o��PP" �Bus�x�4}N�û��'S,����j�_� ��\������o�w��9d�t�ϟ܇�D����K�	�I�zS����]�N�(�s�j�6�fٛ6���,xz4)�+�r�ޡ��X�V��?��~�=��[��f_�L�^�y��q��0��}��. 5\���Еw��5O�(e"��]:
\����ڡ���B��cl���唪C��o��%���~u/=�l���A06��!�u!�[�����s�m�x����}Q���l!˵nT�¯������;�I10ͯ����?F�0�1T���1MP6�Ia\�{�!� ����X�+���������ɀ$����<|��Tю�UO%���( 8WLW��*Z�/;<GG��^X����{/w�]CM� x��6Un����96�;�\ɶ��_���_��qqA��p}�]lo�s?m����!c8@��7�#��a�F�.
1�6�t��*�^]�J�zϟ�8�L6:L���e:77�]��ƶ���]���J_�F��rq%���9_ƅ崋����c!���P��R���h+�	���Z�VW�]���l�d�6	��;>�n��}b�EcTZ�D�y �W���ITls�5���{�
���̋���N��0�%���0g��#c҅&�]����r�U�y��Y�>��l�b��P���3�|,���E���̭'�����zI[�� XI(����O��\�l���`tu� [���Nk��Lxec`k�����Dj�Ƅl�^k8�*b�ꄦ�qUQb֟ ��.'o�iw�dw>�"�4
��8{�7�c��)��4pF1���Ba�����dՖ�Z�;���DV��{��Z-�DH烳�o\/����d
�p���*[�֭d9�(�yl�5�ʵ�'�	���2~�2lj�N%��T����/淬�2��X��/<#SI�Ҋo�xw������?^Y#�G�!�G�}}��CU�ӧo�ۂ�9�̚h׆�{w�?�.Á�u����։lQ�����\<����g�p�(V�c�8q�I�IZY^^�}٭�%$�װ�88'ⵍ��H)J��e���j���t��RlIdǠ��f�[T��ļ�r���c�S��h���T�nN��]��yf1���u���ɩ�w�!p��2�^nnn��! !� ����9����Sv�����A�q��$=W����˳���]��#��s��q�5�\S���u�"�����??1>���l}&�4ޚ��|�t�H�I�
�Unm�3��#s�s�P"����if2x����2�w��r *M宾d�iA��
�=�k�Ξ�d��DYƌ$�s�/�F)0f����=l%Gևs_ ^#����|6��MM��3W��3R�j��~� ��Vy��0��^�5z��~;������M�l�\f��Q�%��t�i�uN?�s!2�ɸ��κ�-�C�ǠCD�$�n�KD������%��ߚ0��x���|	@[w}۲�k��6ZN��̳tCq2� ��%��G.v�On��E�����J���xQ�4 �v���u���e{�o:yם���*�l����W����Q���W �"�����I��R2��.|\__?d'�G~�bVG�t�-�,^�(��(�����imA#�H�m���ha�G[�����}�QK9�N�|�r[�9xEK���"����ŷx|�SΊ�����!�n?�#�;�[~� 80���Fhkiz���S��piy9=�+S+cX}kI}�)-�[!�����C`r$v�b���əO5#��H�/�y|��N{b]#�W��&��!��,��#6sy[�XYeO��d$k��&���U�S�ڥry�22l~��!��A�h��[暖�rX������hX0�h� ��9��It�X���O*���O�b@(zh�H�i���{�7WrjmXe-迾e� dJ�ζʸK��W���R���숒ܚLz�?�[>�'!ܙc��Ԗ���gf9G�����!D�x���G�T�8R�i����bM�p��N���� ($�b�Y��C�˾�)���f+�b�U��>O���5������n�}3������~���ۚ����!NW�/-Unvm�(��Ŷ�g�b0�Z�O���g�'�Ϸ�:�M��2\M�c]�Y���>u��ߌ��݃�̬2tg#�&+%K'.�y��y��i��ѣǎշ�(�����Us?�Yև��>+C~#մ���_��7���&��J�?9�ʑ�L%�S�����z�H��U�3O7p��D��� �S�f��~���~2�b��p$%k�BC��l ��|�7���%��s�x�@A�ה����ro�}��9����''��+
���{��^�W[[��(��jåH��$�|�n�=%KV����j�8Cb��t�y���)��`�1��@��u{�����=|r��sn��E4�~-V�7W'���������2��m�c��8%EEM����+ws��+Y|��8 =�ϙIq+*����no}���NirV/�X����j���Ԯ��|��B���3Q 5559�}���M}O�����x���?�<_)�@TQ�m�Z%d�m�z �x#Î.>�Ǘ�tXÁ�$�������S+o�=��'1�٠�I̲���h��s�K�x��k�wQ*ɒn���S�P��7����-�$�g�JC��Y��`����/M�p$�	��U��M鱅��fv����V��D���u&�ω����
O}��[�6�?4G'*phn��x���۪��R�32x:����G�g����y��Ճ���n��~!{hD2إ.�m�o!���6?���B�U���B3���Z�^�OڽG48k ��`����I�L�}z����J7v�:$�K��,p�aMb�������
���u��������+�)���#<ޒĩ%蟦]������?)~oD͓�����@�w&�ɖ������a�9�Y��� `����2=0������9o��@n���e ���tV�@��B��G�Z�_���[B�^l}����x�9yf�0��q��%����0riU�u��|D�W،�C*�}��˧Ad������#��v���v�#�|c��{�K��Q����V,��/w�;�E�{�wVG�e~,���I{�@ �7F]hHBF�o�@�G��I��<h�L��`ao��+����	��+�>g2�AFhS}��&���d�����K�GJ�v������%�V�L�j;|�l(�Ž;����\���V���q)�@zU� ��޵�=[��{�G�L���[�L1sp�x_f��$w*Mf��/��^��(�9�H�w�Y�(-e��Gr_O�ʍ���Qc0�������;�omVS�_�*)oS�6-���ߥ�Ǉ���Z�r���@�3pG�ưY\R2�-��3����A8�˽�tL'S۬��]�L텐�#��_�:U�Q�\���CIDbڿ��<��q�jˇF~0-�(��/2H���u22�n��L���d�C�s4
���f#�����M��h?�jзW |��aY�Z����G-��� �?tA"'�ϊi񡣕��[����/��`5�h�j�u�b�|���th���&J�(��xz�A�芊���5��7�1{;f����-Ҋ���T��|�nWl�+ǡ�CsM���T��wW�l���z�Y0�����#x�|3�d�H����y�Y���R�ou�sǝ�1�9<��S�<y�����Y��z�z�"� ���a�s ��4M�w_@��<M��wC-�V��8m�W�V�Q��e.�r�t��9p��a���� [)FBpW�S	���H��e�x_�l�H��� n�)VLTR���3���ڝ������AI"]`��8���/4p��<i"�u�t�袍�n~0�H�d\��{�nkG�)�����	�Ť-�Rǝ��m!�?9}r��s�����"e�%���v�ن��@���̏���&;)��e�3ʀ��S+v�X��"ZP��Hs��Ү��6^�����LTB��0�K���.mPm(By;�n��^�}���|����J5V�qz�R��#�t9��B@�])�Ǌ5k&���;+�L䑂�:�#:�� ��̌+M�?�^t�PD�ɟ�-�+�-Ҷ�{G�Q�8�C_�����\ q��X���5�]ށ̎^�3��c~�v>�����}.��aҾ��@ߔx��SBI]�C.6o޽�����`Y*�*
c��M�����ܟ4��bJ�Z�0'Nw��y�e?iF�?�gp����[�Ϩs	�V�r|�/�������埡��ZTS����W�����>�h�;�=4yD�f%��k�hΫ����
���k8���o�M����ghW�\"��fg�U�����!B0�;Ƈ�%��Q���ސS{T��/��$$�% �qx\�WX����j����H�F�O�tw��B�m��Wc�_���x~Ha�D��U�|ct�`��+Z3�v�|
��v	�T������C���U�~�  �
A1[P(<�����9Z�p��N+~��J�Oy!P��.ZxQc"\MW�� HFp��ŋpL~O��ℒ����ާ3LMG�18aٹ�d���\����3�_��s]}��t������Ӊ>����f���ƑϯΖX������;�}Q � a�G�*wC��Z D{��8�ҍ���[m���\'mm��%s����~���!�'��Tq�pPu�_~E�ޫ��7��7���&�r|b�ҪX���D �;�O0zL�oN��ιv{r�2"�9�6�����5g��+Q(��rXȥ�|�wu�5�18@O�Xv���k�_������j��d�s��U8 �.s���I�|{�����΁�	�ܽƥr@��V嶬�\w������-���H�p�ߙ��r�8[�7�E���3�7+qi���Q�E���z�=<J;�jgJ2�/�2Ρ�yZ�:��o��y��}�����G�.R��^��^�`���ʦJ$w�m�`�������i1�<<�V���v��~y'�����b�l\|G�wF�P�p�I�l�"��R��R�����t��*Z��߹/j�<��kb
��vZ���ӣ�"��|y���E��^S�K,�
��o0�l�n9D�zmw�#CK+	�LOZ?������Y�F�s33*|�.�����U��%3p@$n+2��u�*�G���5)�V;ݽ��ֵ�S8�.;_c����b�<� <�����@��@:���W:�oL�>�W#H���.^����� |W�p����� O�����U���{�TZ�@�.�v���N���mX�>R�h5{��CƓ �L-u���Op��w�v�W(>�E��=7��]����f9�y*�V���FǕ�CM�;�&24�<fŇ֒,�	=&`�;�(�����K��Y@� ���\���o�ݟ,Y:�u�LV���P�Ğ_���,,,�p�>&����7K0M�q��K��a��0:����~�	Vr���F�8��:��Ud�֣��� �!��ϋp�E�i�4biQ���S�pb����� ��?J��W��ݻ7׺�}S3j؟�Z��%]]ݥ�eE�/xtH�ukq�X�du��aq_N�qQQ:�H@E� Ą
�����7���P�r����b��b|v׌�ЖY�2<ɏ@x�R�T'���?���+�V���1A�[��V�D,ew��Ѻ�IX6����4�R��ɹ��lF L �������ͅjh�V�lUUUx
@@׼�B�/��1���c�ok[,%)d��Y����W���x�dr߶�/G�^�:���e�O�E���x9��A_y�/��E2������f_��C�K���Q��'!'�)dJ���U iL ������C3o�L�j��S�0��\�`��Y\7�7�q��-�L�mO��V,���7�s�J��L-��Xx�+��;�)�>-'\�󿬺�kS�3P�7F�Z4F��js�bs�B � ��V	@`�%ɲ����`C���*�P��Z���@���k4���E�̬�q������"t�N	��
�<�A�|�$��`$�0;<�vV�&[SG?�ZYm�˅�u�.��j9�c�����Dw��g�˗�$ :�?tb�d��(dU�7�N�n��l��)�'�W�4��6k���<X�����iW2>(����k�s�9�5�7������2J���I���$VU���$ao�\\L ��z��i>�>��jb�2,���Tn��c��k�pf&Dz.歼*���O�W�LN	�H���B��i��,���U�>��o�k���U�~����-���s�ӽ�À*�NkR���Mg-@ӑ������k�X���m�0�ui���a�Q�����I�'$�3qs�\��5��˯����?���+$��kVwE�X]�'�g}���ƨv�IhX/���M�>-l�\>Jr���	{���(�EQ 6 *��HxĬ�퇕z`P,�0�iT�W�A��C#����x�	 �BF�0 �X83���W�;�ɳ��"����2f�Ջ�e�3:"�Ц�~/ ��	BP%��ͤ�E�z�Q.��D�����@�u3�����֕�Y���pt#�%���L 4d�5�;��ǹ�!R����b"{�!j6�r���'����0L{�aS~	�=�p챈cyt���y�S��m1d�co����O���	�mE��~Pŏ�� ���1P�Z�C~�!�Xw�dJh������]v��=��D��D<܉��a�+U���u�dX;�"/�J�Q�F�ηR�S�� @'����˷����!}Mfe�# ��->���m�_�}���-����Ь�
)��y7���Q��:���u��g̀.�#G�i�.�ã��eb����� ��= >�'t>�<,�>S�+<:�4����AQ0�I+�����E@E�� ��?%���ĕ��͙��ϋ�wtǤ0�9TA7\��� 'r�X6���e�f�kq�?����ˑ��o�L�i~�S��<4�"��b�F�3�	1��%m�&M�?��A3�*j�L��a��n�X�N�v��%�%m�/��1&���7��P�H�@N�LN��f�{���>��F�2A(��S�q��-������ ��J�0*�d�ޢ��g9�1��%��g��#�e���	p�!@��K|^�D�{}Exc���*�m$8��ݖ�V3��������?S18��	m9��8�[��(�С?~��D:	������"�Y��hq��G���U���� Ѝ6�++�O�Ő�q���('Ė��|O�/9�V�YO����d�QsҬu��ǜ���se��f�I��I����o�9Jh��>���ᾴ'�����x:���6�+ײ*a��0��v������R
g�y��Q�s��u;%<�=Ie��,f �q��x��F���_a�k�?\�T�K�?�5@�DJA@@JJ�F��<�(��!%�tI+ݍ4H�4HwIw�;�>��Z�Y�{�]�93��'�왯�l��<X�O��������0Ã*��E����s�>�0u��?R,����>�{�����t�2-���E�³�p�â`�%�p�,�w{K�E�xa���i��Q���6�^o�)*k��[������b�����z�������ռ�ypWO"*�r���M0�n�@_�:�͂�[$�B6<XY�����'�����w	�q������b��3@�0Ir����n>��v4�u�=�K*BBx�X?��,���~/��PVi;@�����mX5���[5�%���,�n�s#Ywt}���R�3ƾ�q�-w���+K�Ò�@\Z��UE�?�*��k��jU�����Bª���� /����N���;L�M��vl���w݃q����x�]I���֫c��a5���C����Os�I'.��Z~@�.���뛪������Hĸ��K�d�	���9˿ҭO�r��i��.'�/EiOV�B):�+�{����%N~`�{8Gyi���2�<
;"��{�@������i3�-�	T��ۏ�r��?��[".����V��պ�<���N�\�}���D]=lTv���}��uDgə�,ܥ��?n� �y���/���b�������$<n�M�^��3���AB�M��@���"������u?���fY Z4�S+gp;�wg�ۍ,�����C�\��lrkI�8�o����k��o��=�������Nr�}ᑋ�^5[[�f`P���mlX��������g�@�u>�c�?:���9Z2
�.b�hV��@!���������_W=��@tٷ~)��#78��O�ة� 0C��:zC9ʭ���E%�Dtx�������߻���P�>�Q�����onn�M���.3VN_��\<V����R��l
p8.�:��u��Js�xg������6���I�!4��'�ƹ��fkm� �'��Mw�]i �&�?�N�0�l�}u���n�ߣ�x�Xg�o��]f��[�K��,$U��2~�#F��rШ�>�kB*��X}���(a��%^����)�I�s�i^B����_���P�kwF�;����)�����3[��3tV��v�97'�V+��؁O��Ҽ/�,rN>�TA�nT7&�q-��P3wA8l��w��J~���V���u�  [��v��9n^_��`��P�<0dt�HԀ �6�!�C����=K)�ҭ�����є����V�QK[���'�MA���ӖfL��<�����6��Pi1v���X��<[�2�Q?3����W�X������t}������kL�X�>�v�, tlZ>�W>a%N)Թhu��~Q0&��S¥�&w} ,F"���tmދ�|�s�@�Y�N��ݠPx�;�`��x����"�B������%uy�~�m���Y�D?/d�%;�)��Q(D��'�ͧ�:�?B����.x&U�*�[�b4ߞ
_���3�]�[7���]G�$č��/\�¹zFvSB���L=f&q�'��������P���+; n�3z*�.�H�6��Ȧ	��'}���2D��f�\��6U@�BI���y�3�����%Xt�ZM�m>s;�꨻A��I���t]y])�Gݹ�*��eV{�$?N��#o�9�IUW�C��nC�7�rs�a�i}�� �z7W��J������-�I܍�ʥœ���y5J|۰I8�E����N�Њ(H�~�{�XS�)�%�$dz�a%!k����2��jjN�ew�	��AjR����d��b��F�ۆ�>k#p��\;�C7݀�O��\��H~����Q�ʠ�[����p�`e�!�I���>�nB�e&od�~O�r~��&���ʛ�TB�3/Xo1i;�hwh"��0D@B@�g��T�<Z ���K�����l�6��H/��죮�B��F��C��^;N�x0Za��i�ַQ�	�`M���h�IOg+μ��y�F� ��k3!����2���-��)6 �a�ǃ s|���Xe=��@���pږ���X�@6vo�C)�S{���vvs�<��|g���應G5THHHV��l������*�~����:��:;;��� ���ic���֗���ו�d4]��DM��WTr�a��;l�Q�qlIUx��q�=��xS]-$-���AW��O0{��M�ʚ��ii���\����a'���b��ۢ �>k��fPV���V~��K���0�c��2�Vf����O@��;'��v=j��y+��b��}�g�#���� =9o�R�Ud��|�5RZ�xz�:9��Q��E쾋����:#�jP>~���6�=����`֣��"��_�x���J����S�-+xqq��.��4��܀�$�����=��������V=#��q���g%U��g�	Qۏ�S��%͖�y��ۀ��Z#r�^������/RRRv �����!�~#=P�����#:X�FTƟ��e�l�.�[�]/���� ��
���W�:�/���m�ԦsC�|�н�ZX�������J�(�Z��k^��g���������t���+`!)����f�C*??ً��.�q|�>�qT˿}����S򇯷qe'|�g>�R��e�2�M7{�<�?�X�)900�Ǚ�a8P�=<Gijz��.:��=������+��?=<�cb�I.%�e%.��%�8��Z���p�N���سw2�OfV�lMԨI6���i��3G�ʦ�@�d����g��N����A�~��T�|�Է�2\������c�._��%���ѣG�蟚o���s�����wQQ_PSJ����Sj��~ᴦ���ÑF�- p|�o�/�q�5@u�g����N=���޽K�X:���	����^+�ƸQ�\��Y�n�������~YYR��]]��v�����r�h�F�V���Ρ�]]�&V�����
�>��4�M$��HII����JYP�aN�#[�sc]�h�CB> B�622���q���E���&�fLL����ΊtT�����3v��߮m:�~}�����=pJ��3u:���95𝜜���|��t�ҭw���E_>�66A�����9K:��,��c��o-,`E��C�h�ݫ8��h"RR¢���\:���������e���획���9�=�� E�1=f���"�Y?h�*��< ��ܔ��;wHiiŇ��o�RW�G��>-M��ull�������C+�MF��-��؅��q$/�雁����+��C@�nr>Oru?q�,m�Ŭ��	==��43)ٮ���ވ���L�~�B��m�]
������W*��8rl\�7&''c�վ��ǯ++G�=Z�������8ՠǜ���Mz%�rrP����[TO��H�`���ݻ�DD�]1��(((U5��X���敼k�����z2x��������S�3�dj���^���	����P.��="���ݗ2VVŽ�����
����ӑ|1�޼ie���o���~�~钚��꘹f��{����=|ghI.�(  R�ߕ��((x''�	
��n
�{��j6p�5��%��c�R�>S�0F��e�E����~)�s����qO�������^��t���t¢	���OD��VX��ڥ;������n�����/��N���U�ժ�S�ⱐrǯ_QU�"��d��Fh�!;/c�#0�^�}��g����5!�͉;饥,��F����UԴ�M@K��F��l	$�٬�2�zui؟**"!5=4��m[s8\OK�8�Q���T|��Q�3P�ެ��o;"�bb���V��$#�{5<Y�%�qy��Wcc����I�x˛��_�z������2��+a�-C��HI_E"�c����n��B~�K�&༊Y��XR�o�\�$�1�����z�|h���$#/������f�F.��;r
�ssт�N3{]88 <n!+h9����E�Y{�w�1Q��>�R��"+++")����^�-��������&������O�݅vE[[ ;j�M�����ϲ�bd�TVVf��4�ݤU���9Y��pFP2�p�H'	���aV��5���SaC�
�c�WH�?*�$@��.�]^	Ivwt�ݖ�E����g���v��K�^�6~VS��Dk�����Z�/Fܵ�r8�ns)��g�g��K�VP���/*�
�ٽ������U[[� T��jFR���A���#m�5s;�F�''�.��i����u�Bh^3�h}� d��d�_K��j�ӧO�_�ĕrp�wg��p+ji6��#�'`Ƣz<%����N����)O�'m�KM�J��1-n�tt�|��\ �իW¸Zzz���]���C�����SR^G��H�sx C�-�wl2Z,��^Z��X��������0pD��Ӣ�ޚ?o�o�YY�R>Nq��6���ť8ha:I���������ْ����`����w�ȃ�&}�g�)4H��w���L��
��|t�9ź]��q0\+��
��k1��Qs��2�|y��]���䑑�t ��iwq1���B���@#ql�*�t�f��H��h&J�!��"���.0j���H.�o��@AEE�Ʀ��c�Z����G�PQy���Y�����o�����3�^BQU�',,�9@DÓ���G, >����v��n��5Q*E"����d���g�����O�j�3@�Y�x��~�u�WȧɓiN���;y������9k1S^A�w���[��a��l��H$d���2��uT�?�Z/u����R�r�����.�uzw��:��W2����x&a}v��Ǉ�rλ�f�D?��\�=���er��P{����?�ͧ �B��0�z@Hw�D;͍�	��2�S��Z6��̣�6h%(���&��6D��L��̜g�ؘ�OXx�n����Y	���e�j\-�A097��l�Ez<u�_�~�6�C��u�P�.V�V]R��^IN���e�0�CJ\�ׯD�U�̔>ꚓ}�&��zرY?���o�"gf�����orr����M���]���=�^ɣo߾�lm� ��%���1�U�mmw==N��#�tު�X�
�3+'<9����gA���� �Ϗ��êwv�W��˿:;����u���@aҭ<Ѥ����**~��"��n:�]u�ŷ�%��ۑ���N�%@ �,���D^B�ћf�|�yFD� �.��F_mjjtגW>�=;��|�q�Hʴi����XjBF�PpHH�e=PP�F��^�Ө�]�6[p��*�7]�=��z���5w�8���1�g���#]���C�"���	͚j���mY!���"��+9����,=�@|��>��#Q��线"[���E������qWGH���|Q,-`S6,�e��X�5-��+���tt-�^ )݂�J`�;;/�-��+(������a����V�䥣|u=P����D�z���4ᴖ�����11���}E*��p�>�1���677g��
�ۗ�R��3��G�yrv��>6,�v����-���yjT�6�Zpp�?F3<1Z7q�p@SՒ}��){�����Z�O�PU`_��Pj�X}0	�9,�N�����h
�����9.h�� ����{�n'a�.S�},�o�X��l����spd��o^��!""ʓ�H��/H_���3��l惎N�4;�&f'��	@�>�2{��++Y���f���.���{�~6a�^Nr'&q;&��gcgw�h͍u����k]�&�9Mwm�˴��b�8XDӢ��顤���ـA-ӝQ��Q���������9�=X�נ�g���V����+�JL�a��}����%���������=������LLɆ���G ���o��s�𲭭m��e��<�e���	nn+����u/u����$�*f�т_��Ztb�ۯ.��i��z����N���`��)=+��	��aIR�Q�ѥ�����!c�CB��+<Кg(��ۛ��TP�ThA�n�g�ffe�t�PԱ�y��#�$$�'{��#̣�Tk�XY�����*r,��C����������/�����P�V�"�7E���̡�!q��k8�igϴ���B�eӖAE����RS��&X��wW"��������G~��l"�9��EF�,����F���W[���OY̩N�'�E����+�Uݹ�TU���������%����:+��/��!��F�ꬩ
x����&+�8�[ﵢ"�R�ʷ���濾�i:k1+?��*eTT2GO���_'�7�\���xz,%��\A�K���Zi�y����TXw��*·f�������ARβ���󋰰݄��'��O�C�#�yh��i��n���v-�v-?B�~���%�<�#�s�2�9��4��?� X+���y�{e��+!g1�hU�����P��}B����y�d����Pr!�1�냉6&e�4�
_`V��q�oM�Ʋ}���	??��I�2KgE������,���B��k4�6����),�,$<����~�\�q�U4J����d��l�6��`b_�IwRNv��&7x�ګ���៵��J�ws�m(Wbe|'?�	&"]
~�P��f/�Vd�h������ޘA�ݿ�3t�|�����W|��*=IIt��)b�Y�,��o,��5�{�=�H��L9�1���E��}�LA��^ܫ���/�"���r&&�6��F�(\���h�)ng��+(eq�+,�����[�����H����H���e���7p~�la��v����}jN��N�=U����v�W������|e�N/��G���IO��C��3�(��h����������5Iq�X��ר�v!�$��#V�|rv�>c K�B�T��� H���~��0?/�h`$2"�	9��t�on���ƾ�[�dQ�.P�@ ����p�q�]��������6��U�_�Ar�<m�A �T�>6������`�·�[�������;\��-a�F	���3�0�//.��������* �£N��;��ÄN)�~� K~����4���YZi��H3VV`ҥ~�����3�欬,��ٜ�|X�~��뗞������ޞn�����E�m��V�m�3i�c��i�P�Ӏ���I�;����	?V�%��|��J��wb���w��J$=77}5N��	&&�:Ъ�$�HK�����il�vab���E��~"�bT�w�4�+Z9T�MA��L�FN�j�v �o@������iT)��+�6���5o|C�ѱ��?`��.�ɴ���no[��E�p�]7l�\��f�w@TTTR�k|�,B&�Ac��VAFE��_hb�ϣ��Yk����jq���r�o��8��yͻ<d�ˈ��1�����2���;de���4TǱ�����D���]���n�GDD(������pĐ�zh����TvK�ϒ#Z�U�8u��oۡ4���vʭQ�d>[�<r*
33u�h���X8�����ZZ�`$�E�����G�)m�g����� ��e�q���&�ҾS��[�OP�����iqQQ�0y5���^'���z����p�Y+n�����R?l0x(�H8Q����s�x����
��,,R�{�������|�N��FUDm� ��.7O��1 ����n���]��'E�&���2M�>�**R�D/��:����Q���j�^�����������nt������!):��������.��u�j����De���;7C�7A
5����i�m�П&��d�gKqt�[{�RI|y\L��	\w ��kW��XYY�D�|���!#�=�?jFF鱞����-� <~LSU���^��V@	u��q��,F=x���%���5иJXV�-a<�8"2�$If��mHG���/�M���G2D�f-�/X��ڇ͆���)m
O�MB��=�Z2�YͼV� ���W�i��:�f_�2d.pi��O*�ճ����*��j�-aa�!<a=v)_��D�?*�1���E�l
Vʈ�ʆ�	��f�-9#	��VII�0橔b�@��m�$~�� �2�I���1���!���%��2����/��V<��ͬf$Ei ��<=X����r4�a�V��^�T�3���&���.�# 򆣂u?�w�02b�[�t�<��ɷnNL��U �tt���ڊv9�����M��!=�4*�79��w�`ջsѳ]������;QAІ�R_��ƭ�§�&/5-�]���<5U�YL���2����[f�t��")}~$�3�_����ZL����X�������<��qpp��l���@@۫c���n��aT \�P�7]N�{H�j42����T^-����d��!C�$��o�J��<���S4�`��s�<G$��7=��~+�����2BBC��i3ı�����L�]����"<46�ނtDkYE�8i�FH�d�^��L;1_���}���Q������Lo�ǋ�r��Q|��z�`��)q�O��P�2���k��¿���i��N�T��r�K�'HJ�2�x���0�o[R���w;�yq�n~<uT�K����4~���$���?��;����G�x�({t��Ü� �{Xx8y��/�R��I�2"L��\�A��+C�F��	"���ïm���bd�Un)�N�Y<��oe���C��|��I1s��t��S�6-�xc�8]�P�(:Uύ���Q�������>qA��	�]�Ȝ�+z��^�
��b������ǜ N��}�Xk��o�p*�/`[GF������#�$�UL����u0�[#c<~il���u�tR�m�+�c�&���5L�}N]g��ß�Zރ<�+�]�>��f�STV�pt=;lX�!��P�	�g '�e^wB\���*t�����IT�2 	r>>b�iW�x)*X�Ȑ��a�p=evnւcƆ����~�����&3�!�c$4x�`?�t(���@������U�HdRR�'��&j^�	��KiMM���->>jҤF�*���KJ�ÿnM��%5��N���=8A(,�ݹ���	>��br>
6%5��$g;(�?�HFC#*�-'.�j�7g9PP�:�fWU����j�		�.��������C��.CFשÄ�IF�q�}���·�r��`�hi�m%c�'Fg�j���{~4�ht�'������-���j�A����X;�8!���Yҫ�~c/g�9V@N64��0X4�+�gѳ�*�H���}h05�qCUU���͍��,��Jv�lp�g��6�> Ŏխ[�����J�{f-���<�~Q�^�	0�^�1:���+���T]��Y(k�'CT�s�kNĹ{��Y-gbAU����00�������wZ�=޾J2$76�`h8;'絴t�v2>=����ײ2Ł���ĵy�b��da�z%���|}:��_��b���?6D���$VV��0����q���<"*).�����cxq�n����O���¢��JF�(���a�;<X���Gx9�	J��B͸��A�Υ�ԥ�F<^�޶�uc�p^�����}3N���HLD�%�ZK�MMM@(��3���kəv猖b��nk���3���v(���s;��(�aeЗ4�rq!�5AT6�/k��"���a{8�������*ۜR�#f�__���A�ڮ)͎
�`���k��|���j��S=i���(�N�	֟���895����`w��� �k� �C𒫁��S��xRA7�4f���e.9y"6$b<a�����Ɩ3s��;��Va4�F�M�S%��ۓ�]��3���uL3���4%���wܐ�8�c?�%&拥�����"�@�����蠙��+RRx���K�qi�#��_KJ��*mcJ��@Aӌ":����+R�m�0X��E[yVʊ��OϢ����'��!g�g��)�vCu ,@v�s%ܨn��]�k7���hݎ��y1Ry��l���=�͝��+���p��r��������\�����!��2����U���eQ_��-	��RV��\YMMM�����Kh�i�J��DG1�8NRPP��zzzj7!�V">G[u ����N�}
i1� ��H�ڗ-����oq�����999��幹ᶌ���s���<�����돦�1�;{�x���b�����ksa�
�����O�K�;'m$�ʞ��R �N[�
�M_Pq]��V�I�D�Z]}���ab����(1;;���	���IS@c3���tx���O��U[�3�4�-�Z3��U���!G���Z\��1>>>jLn�ͪ�ϖ��N�Q6O[�����,ZͲן�����F��yOt=TE��4N���ul�U��C|'>Q�"2\+��#$!	��^_]@D��p�-�V�@���؝�I�&Rffy��(���II[�I^v�4���ayw>5{����8A�wӏ�y�>A� ���>����hm�'O���-�����߿���fP|،�t��l"��h?JA~�v�kkk׹r#�����gf�h����\��=|�+LUK��>Kg}�B{x�"���(��|.*bvJJQ���-��FM�E���.p`��::v�<��m@s͟�t� �(�N�M%u�Ҏ��}|@Grv���&�P�[n�cSe�%��u{��e��߹��KY�2#��?Y� �%5�)����ml>�̵@B�F�v�d���-H�d�}CC>@c��!;�++��[S���L������ͪ7�hF/�PQ�۬�]�a�_��jj[��Mw{{(�%��ﲻy�����	)�d���-�.	����i�6�/��	�B�wGP6�)%d��4s��T��K~�4u~x��o�P�3-&2�f���䛓� ����"q��K�d�����n�b���|�\�����AMM
�u�i��||��PFZF�7ZZI�!!�s�ʥ�ǀ��b���B�C[��&J�8	J�߅�u+�K�2Dv�<�[/�]�� ���^�N�:C׋~mI�;%�ë$#[���caO�������#��y P�f���I3|;��.Cէ@�t��@�Z�`W�3�K�R������-����������m�,*<�Q�������.��mljJz�����G���$!���
JJ r���f�Z-��� Ү��K�z��m�4@hX�w�)]9��R�==�QEEE��%-��t��Z�%GC��O$��;��������h�����ʨ� ���JLF�߼Am's�����IG
����O#*c�_��$��/����Zt-,�;m6w2��g�YhE5ВMM�޿O)=���������t+���'w
`���F�wE*�R&�:;ã6�c1D��H����O̡������9^GQ���;,�E�R��!ѥ�<\��H?�/���l�J,#r�诣m���n�ߊ���U!�UU\��`���dX�u#��.4�O�΀�����J�m�����^�x�? | eunN��`�F�����e��[�<��*++�L��f�0S�Z[[��Oq��M|��$���I���l���ǻ���ù�TT�D��u�8;o?��\������nR �0��IRG��Ё�o�F�l�}T���$ʍުW�B��
kmmM~�Iu�É��z>P �з昗�"V3&\5�C��F����� ���<|��g�뙷D��K�[W��f�j{t���؍v�Z�^�H|����|�����P{? ��\�//�#��{�n, ޷O���{�����p]&p?���g�W�|����"�ۤ0߆ � ;�к܍�Z{n����6充��;s͍�#Z�#����s�wt�E%DG/�'��)�nV�c�}͐����	?��N� �@�mydh��G*g(@�J@�� "�o}Z�N~~��Cȗ�6��T�w��*�B��q�s���;� �&��5qX�����)��99��޿�V�#�ʒSR�	s��98`�Q,�]A�y׵�r�g�w���f}�u`]Yq<b���7Β��@Oy������x�h���u:�*:�tz 5 rz���&��ya�����p�M��a���3�o[�\N�_�:::���m�;:꿹iVZ<O��6�%'9��]��������Ԍr~~-�|9�	�[x�װ)�ǧ������/��6�$cv�������-�$l��>g���ǉzE*�nN.���֑�|�U����c.`:�#��?�:=�ZF>o�TV8ѝ�a�57��&&��R�W"J���!�F�Ɩ���<�{���	&v��]Łί�%��?/L�����J(�&�'!��(A)��f�ⓦ1����%ť3���}pwƎ&)�ϕ+]:ɭ�@�a歎�m`�,�'-8�]�!��ռ`b�<?w��l%j,/������c� [S�"�� d���r�,ⷤ��.�����n���&ͨ�u��f�v��@�V"��:#q���Ru����#�,F �� �
VN�Y���^$l����Z!����2+�m[���X{�DE_��<���g����F���t��O��?	NAռ6v
�4Q�~OT�J`a�s�)o�0
vv|�x>�I������[ ��V9����sul^FU�>G�@w���A����A��f��Q��;_���z5����T�#��qa��S���Bm�R�k	�W��B� ��dW�����*O��v�Q<J��Bӊ�������~��k�P����fbb��9A���HV��ӣ?������X�w�ӆD����}�b��j�q�r~m�|44"�%��Dۉ�qi������ȹ(�\���M�Q�yg��~��{<nC&}}�����q�*�􆘽Tr-zd�HM*G�G��a�o-�jfH����F$�)�G?����>���HGi����h%��^�m�훚bxJ����ZrS$�^��D��S���c��:�o��!/��ृ�ǯ&$<��¾�#z ] �u�qĀ�K]�`1f��o�JQ0��4@�'�_j�V �pه�ɜ���'�w��VP/..4 c�%1�T�෺��qs�݁���	����X�7
��������G��4�/^�P)�����gB�~*Ě��$��+,�U6����5�0�i j�uO:��/�Z����vV7Z@𽂪*��:X�Q-v�/��7o�+'X�� � c�n�SQ��S�!���u�#���ˊa�9#,,��F���N6*P���
5E��_~ji/�D�ؠ6[.?���_�X/��7������&����k��z3(�1ف@/>3q�a�������!l �U�RG383��-N��K�.{����=�W<�ǭ�V��B1A�i����\\\��P�(/�R+�V�ǟ�۫�6rr޽��stx��'�W��l��RFF�	�Yz�YX�z�3�ֶLVH.V��>5�,͕c�Ȳ܈y�E]���	Z&��SL��?�����

!x�i�� �Sc����Fb?�J��M�kiY-��ˬ.`��{�@r�>pxX��S�Rx��s��S i�N+�.��T`Xŝ���`l^�x���.?[[Q{�h�۟�Vٙ�嗚���V�!���^v"p����[�Z
�;t%p+;l�<
6���E������ׂ5&#�
kO���3�����;��d����I���������(622�^P74�
�L�}Nh��޽~��t��u��~���t7��/[.lH0p1a�+�.�^g����F��թ���/?��=P$Ä��-m���X��ئJjj�&&91;i��R~�2G⬌�+��㩢�����M���B�+7�/$��D��(m��r��NN2��00�3Z>�t7� ��@cr0�K6���@�EA	�X�9{���.FzzI%`ss�Ro�=���q:Y�ہ�:[��ĺ.�>'�KO�x�BP�����1!!��7���ad}ۦa���p���n���9>�(3??	X6�����<��gS��Z�Ĵ��?�(�ml�9e�vvwG��ą�z�O9�Gw?e����ۻ���	`��F��T����[ɀ��i������QpQІn���~��9����V���ur��`���e �=��9eX �U6ﰰ��Ԏ&vOϳ�/ɒ���<����#9+KTd��������Sz�g�#��ã@����
J�s`����Q���&�Ʈ�F
}j�'<�B�j��qTH|8���v�]v�����5���ź��@�DHd���BxP �ڳ�>"?�GKn���������~��X��xx�r�S23E6@^�=�]�+�%Ƽw�^��q�Yy
hk�y؉	��i�H�1�2KKb�x�W�+��66�������4��w�?�����A&#���m�����
P^�k4?26�)���Mop�	���ί�W 1&PL@@��b,$*�_��Cl��ĔlE�����~�5+lt)�H���n{,�yb��<` P-`۴�Z����Ϗ�AQ �U��2��@C{��a�ld�'��L��fl���x/������uC8�쏐�S=��D�C«�啕���<D�r�6cY�mX5pn��#�n�~n�})$�aZ��!�������Ma!�Ģ��S��|o��q8l]gbi��/�`漣Ғ��'�O���3o��y@��Z���(X�q���HR]��R��^�4��^G�@V�bg��-�qMll�͞zh��iia�T���r^}�&&��<��Z�6�R�Teee尘�16>��[�Fpyqq�a�
�G�� K�W<ϑ�-X�]\3�-A��H�����69BV�_Ua��ׯ_��
��ePPR�#��ob ^Y.���Z�\=1��7P�!7�;::d���Ѻ�J��N�w�d/�?8�i�%���q����3k撘xV�5�W�`�^���3����4��H�~]��{���ťs�0���C�X��d3ɚ�Bm�K�KL�`��)X����3"b��W?�lc�����������num���_nЫ}i'�40���Q赆�<�`A�}A�I�!Iq���4����=�C��|*����A"[`^��zMV�Ӻ9���!y��+�[}~:<԰�0o[{���2E�a�Ȉ���=�������r�4P�^��s���)I9�	����,tq�C�D���N�[�����%�N6X��۴��3�|�;"imY������DSS�x���[a�ꕇ�0�;3nK=I�<�,�=��\�3b��E�F~_7���Ƚl�0E�.�3 ��@ �$�=�?� �Q���̗����4���g��=����*5��6�NNN�ςCJz���2@�O))���eY�L�F'&����	0������/Ʌϰ�¤BWr��'���xK��z#33�(�I��t��gar��J�3kqי&x����b��z<{���(�����s����\D����bcS��{K����S�&��]+ȟ�_ڎnE��k��P�,θ����;��њ�ݰ�i�J������W��bBFF@�FU2p۞�L�򺋌�>���-EEm�{���_^���/4����}tW-Ê;a3آ�39,Ǫܺ�$�Z����L��YpS��� �P�Q01[Ƀy��������ݼ	�*^�hZZM'̈<��`�>���i ��5�F
���R\�SanpK�A�@o���u66��f�����8��f���寮.�Q��0eeߠ �Q��ӳ2�Ī�0�B��Єf���o})�Г��[���OȒ���f�j��#4׈>���ɞd(c�@�iW|`.���?�����o��$S��I���!��]�kv�߷)�k��W��m{�85�pq�>ܬ�r�O�F������5Ë�`��5�����e�
�^���~C����tV/F��2���T,�)|�o1N��d�'�=���eb��T�}�xxb�v�v�u}y��a��CC���^Fﳌ��[���a����=���z P��{K��_gon5iC�o�������:i�*�Zr�'�RT Q|��������֋k���,���{(((~ ?�`uHR�).���B�]����9#���$R��#��`����\��|B||_Xゖ���_AC-�o[%������䖛/�V6PxQμ�)X ���&�E>.**j,�����|t�$���?ee�N�h��jf�B*K*�?δS%�(/�}Xk���e@�?���6Y���9cGgg�N�I�:`����T��;�@*�����O�Q�?�^vb]\^��+/W�wu�����n��?�m����W7
{�_�i�9_�+p�t�����7䔔H@��$kll|[�r'���J��,������geaE�íⱑ:ʧ����9�঍Jw$���+F E��03V��J����Ùbb� Hbz�&�220�L�O��1rp<��9(2gN��ǐ��405=8�1��|��)(D٧�a���3+���{����9>��(��:���:�7A�_��^d�G����};-�Ƞ�L[���Z��4�aȈ�~ E��b�e��X��iw~ #E�[1�y�T@"��\�4�;��|����Gy��)<cP,N�l���-$,�q{��K���p\.��3��=Y�W���� �a5��}���H�"��M1Of���`	�R���::3���L�l�g9,�)N_��
�?==ũ��9��"� �$�|�Z0�ِ�Tg���))�wx��P��`SJ��鏍�<K>���Q֎���������V���
��[��U�:�i�.��152�H������9�-mmwjj}cc�|���~yyٓ������� A���p�>>�򅨵%l�x�]�⽄t�)���4q0�������+�`<����ͦ�4+��{��,8f*M�x6�=��6��	[��,,8�����9��V33�5x��)k0�C#��M	��bRN��65g��NW��7��Q���MK;I &fº�W�>̐����.܁fϧ����DB������2yd1�]z�J�*j浸{K��Q�E�����x{�oޣ�y����uG�O>���Ϗ��xԀ�����}tw��xN����[%pt�Hdo*P�Ru:��?� F@�=TRR��R�G�-iB�>`��c�_�����ݟp�[��V39�$d?��j�Ǐo�OK�pR7��\@3�%ߚ0�8�i���Z@�΀I�?��j�e��KJ�:?��������������׍f}��ѮxN��la|o ��M&������y"��!�\FDd�{���Y6�C�nݺ���ްQ>��3n�B���`�E�:���s����QQx�M������]��_�G��H�'44�c6è�PQӖn���WK=��n��O�F������߳�p�T2�zW�G�Km���y�gF:B'd�N<��DGG707���Or�Lkp�+;���,�_m\pxDo��ͨSxt���V������w��3�յ�Y�?g1�	�${z��fO�3R���㟀faay��hy<�uM��.A����ߣ�_�$%q�O~x�Ⳍ��T�tt�620�E��7�O0ax>�ū���bt3����� '��W��Fh\'#��>q�u�kt���>���Pq7W����7W�C�ƙ�'������b����X���{w��?~\S["�p���Jv�h��P�22�أiS��;B�	��JV���۱�1���^G�������������y����|<^�i_��ߣ��f��3\��;9�(��R���q
K���w\k�Q �w����5@�5��O��G���@���Ǜ�@�}Ψgᭊ���epa�⻒��3g��>ž�0�_ҿ����u&��)b�����
��7�ô:����>������ʲ��w�7�s�ە+�NC7��g�� ,�Ӏw۳6$*�
gz~��F�9�4�ߵ�&F�O�XWCçצL����A�C �T9�.�u'>���K� �W�0z��i��N��Nܼy�OQ�==�x%�[���G�����vsfB�����*��KiO<�v[M-��P^�ŋմ���QP$Ŋ�ˀ[��/bb.��#�����m��F�Gɛ��Q�;��x�wr�x0�ș�����L��D f+�tz����[JՅ�*΃��n#mF��
���������x�@IɁ���'E��}��3'
h0@�"�����K9��5�y�?�e
�,�����2T�/M|c��_P�����:�[)/���$ޡ�?v��u`���^�8�Yi�"]�2����0+yec&���5��Uq�߭ZE�y���0 VVW�7S#��F	X���ba��C�Ǉذ

��_�Z0o~������J���e��=��7��oAף�]V�ஐ<�����Ks�htcڥy���%���4w�~�=���:ImP��	b��
��-�ʅ��D����i�E}N�U�;ser6x o�h�I�L�<%+�0�3*�����$�����>�{�e�%lI<���Yȥ?��@'�q����CEEE�QՉ�[�n���Y,�R,�N��xy-���`x�U<o����5$J�h:}�dEڃt���%)�������Aq�a��W���;��p�ѡ�.��o�̫���,��Ÿ���|��M@��r�Ν#GII_�9;� <8?==͟!���]�5WD�N�Qsbc�"</K$�*�*���p����쑗 צB�vt��y��:�<��A�s��Y$�W4`g��Vꡂ(U3M1�cU�Ց�_��::� ��i%�|Ͷ��@��A��^k@�p���Lǜ��;1To��g7 #r��8BN~3�{t�jy�#��F�lZ/N�I&�@��=\0hx�X)��T@�X�/#�7^�S�pummN�ӊ) L�/]�v�@0�f{���k�̸���s:"|��Y�W�G������\�R~B#��æ�䴅PT	�p��7�233�GlE����B"��wo'%%ŗ�S���oMQ��њ7fiiy��8q�<Kk�̌s�����ޅ���>��PQ��ZO�+��W�����[�Kvz��������8,�S�0����0�FFNN��\~�n5���]F�[�&$$�^|����
#�e�G�B���e�IIGlJ7�_����:�r�3f��&�xL�����r⁈!2O�[�Z��
�{jj,E�e��
��<i�wj��̇O$�~ ���\����=y���ӓ�����L�������jk߆���������W����" ��]/�7;P����-���$�����XiJ��!�k�LKG�lY�}>���yY�)��y�֝�G_��u��+��+kk'�U��;[�Ϭ"�tJ3���7��j̗����y4賢�?�����G&gf���5��������5�<Z���E�i/�-���x�(�9q��DHHH�u])`�S/�z�X![ۇ�c�g	e���y��χ��o��*+�;�TY)	�24OD��[x�0�Kb.�e�Qo�R�]���U���А!�/�/���䇳��U7^?�]60���KrzN��QX������{{��EE]4Դ�/��*q-�\|Y.�4ƻ׼ �q�23�?_y�,JE���l�����I�N��v����1*�3 ��c�q�Z��~�6������w�-�,����j5P�+Dv�8���$�U��˞C��\����;����
���
H	z�i����]}9��g�3�v�RlT��^$'T�׏O��>w���<, \��	�^щ`� ?��@popͧ��~?������J�~�WN���)����B?�������h7ңG������̲5���t <���쾅�+aH���L@J��ExE�]b��c�����9��	�4tx���׍�x7�B0Q���>�JS��U�����p�d�4s�������D�/k7�;8!�^MXw}��O����6=�u� �nS^���[Y�e]+�]I� �����>>g��&;s&���������p�D��`tIف��I��, �@c�s�Իk7�H���#l��c��X�N�ׯ�-�A@��[D��v .>a��?kzX����w��)��h�ÈD���U�g`��(���Ł��Q�E_�.���(�3�d7��@ò[7��@�1����>}z��x��ъO)5~�ZZօ�2^,��k9Tԁ^�� ULV����{38h 7��rsr��̏�sq��߶uɷ��R��1���b���xv���QŻ�#���W�q;����[����'��49��;�<{�{�����������:T
|] �5Cg`�RZZQ��e'Q'�n17~G�SU	q����[k������N��Wo<�s���_N��-��vvv�!��m%趽XC\
��P2(u���e��>V�$�x��ϯ��Sr ��$�ϒ���ů�ɘs����qל,Z�s�c�T��2�G$���bp�`�:0-ӱⴐ��i��A	}E@���a�Hw���}x��4���Ov/��ׯ�PN=�j�K.�������]J�5�U�s@ϟ��l^N����@b��p�X�3�4�G N\��?"##�}i۰��Ύ7�q/'�� c�ǯ� ^+O�@�86]=ѕm�wcs=������*�~�vu��Š����U����.��*�A��>����b�)���u��S]-ϐ��=� !�`<�g<z}~k�`^�׭�6�mڨ*��3�J._�7�U�9�~����胧[��k��~�赓&��?�|g��ן�E���a�'4��wl�ə?>Z3��$0��s;N�Ol�}�.��qh��9q��Y�	�8�;�?C���(��+Y��L=1�T�\<�_��s�f&���-����[l=��#�;%e�������2�#����ܤ�K9��A�Trn{�T������0a���&3�6�g7R݂��\�l�����P�sss	s\�Q��b���F��|�	�N~��ܖ��g�";5�r!�=�HEs4Z5��<�(����4��6J)ݚ�ߎx!a�G���wN�[O�b8��g8�0�,&�J!���"䬟����#�q�7�V�jKO�$���
K ��換5I5���&�=�a���
��
b.TP���(��0)A�t�ۧ��N&�JT�9 ^/Hɢ0'o�M��0�h������G�[����%B�V]g-;2�FY.%zś��0�zW��'T4�]
B}�{�5��p��R�Q�l�w!�t�3Clp×&���{����-�]ى_r՟롨����W�Cf�]s<|6:W�pq[El��8)�D��@�2O%L}�I7�T����J�x�9�ð�Aq>�PՐ�z��h��φ���N����R���+�!�>z����5�dU�R���<z��r���Ũ$�r%����s���k0�|kz}�U�����Us8���?���n��5h=3e�������	�E}�koG%�\18���v�N]G]�"�v7|g[��Z>����ZPXX(��0F���b�09�b��Ѐ_��WF�
��~|b�>(�&]˳줲'���:���imtV�o4x�j�b�'b_�<Hvy@������M����C���ש��o�K��q�sa�0����l���῍qb�0A��bz��y���Kn�)_��;94}�O^=ejfv�-]�{�Q�>�/[�<=���������u���ى2^L~`�Վ�׆O}��.�J�Bu[Uǉ�ʊ�&E��rғ����]C��'�/!��r�PꠝIIN���q�,s����İ�_V�_IMM�(qYmj�!%!��0�3�8R4�c�ͫC
�dW��-Q.���&��	����Q�>�*��(���o�wHuuu�J:���J0�[U�O=�����Gp�g�s��H�:��a~�g|�GEp�|��l{�T� Xqjݖ��ۍ,,�X�i�+)��'ZP�:�����K���c��2;�<m
z��yx��$�=o�۔�v�R�JR���V��V�z���y���X*�c�g�u�o/�T��r����x�ncy6^�����*膭���||�_v ��&�Q5:�0 0P7n![J��7�t�@�'E}�:��SO�x�lo�qrr�sE�Q0��e�)=~z�a`�pL�]��ė#�P~N���� ���ts��uN �M����d�t���Yv�Z�~a5[mS���'U&�����w��"~kd�צ���-¢u@���S�\*���#�)��v�����k��Ӟ��Q�\6�ҋ�ذ0�,�`M9�q?P�B�夠��^O�|Y7	��?�-���6�o5e���W��o�Y�ڡQ�I�}���9�"'�z�'�����OA����*P!Zp,����T�l�H�=|��X�Jje8�����fGN� �X�
L�N�ȅֿH/9�L"�z�F|SZׅp(�3S��yx7��7.�L����疔$[л�2�;��V`���qP�lt� ?l���Mb�*�>�����,��_~n���\�na�\����D�U�q�F�9,K�t^��]5���Qg��|�N���/�	ص�f��?�<0��L¾�IZ�/J݃��+A���0w�mW�����J��J�b��	�2��wK���d��4K;(�8���X1N����3�CY�EHM%[�C��h���%���<�ȡ��}9�>a�Ϧ��*��KL���cϊ���b�dA�&����o���bu�� ƛ��tt�V�C����;�Ď.ᕈ��[i#�GƲ#K�f�|7�"�LIѻ\��Jr"�"B���u;�s')��|��m������k��-��a:�tU۔��
zB'wӠ��9>w���V.�(v�|24!�>�"�cg�r��"�8�I߱�-���a�z*����'�w��(izgf0x�=qnK�:,�s��� ��� ڿ~�{��k���9�h���J��^x{�/�г;]��c��"
)��C����ߡ�÷ 97Wa��#f����|q.ө�4�©�)z��&{����K�
�U�J|�9A_\ �@�����jy�aG4����S�a&�ƻi֎J��_��Ѷ)��������8�6�_����ɳ��bތj�P5d|xt7��\p�X�U�T�iS�΃�Q�tH�@��<��")F,9ӥ\' �Y��8�m�!Z�(y���8֏�E��9'�BCC#;\m^�(�G�`\��互�E}ܳ3�+�I���g*f���ޤ[`ݗ�B�~%첂kS��l�棹V%�J�D���xc'�,׬���s��{d!0YC��.@��h!�7�u�q�h��x�0kS��O�}��5Rh��?�asqǋ��3�� �#rmsO�$Œ?�vd��pi7�P0��z�\|ra�2�p���݅f��@���/���-��q���|�u��/k�،�z��y�B�a��V���o�_ YD	���	a^>�@�1tbG��߶�ڐ�k6j�R����Z����~cbx�6��c-������l��p���|?��״0S��qK*���%�����o���ڙ�β���mߒKd'|k:)H��j��WI^����ڀ��#�_�;Z����s/�m�e+I<w�{�K�W��0����T3nMVP�َ�v���y���eS�����+Sr�_�'P�[�̍f	�(��z녝Eə�E�ℍ&���t�RL��T���_w{a�]uI^5Q��/qy
�IO0��#Rv�h�Z���=�{u�On>rr�G1Eu�n�>����b�jޚ���6>�0H�m�JX�Є�Rh| b=���^#A��ps����*\&��@i�˞vY�`ѥ���g�s�7�Q���Ű�q�N�������޿�{� ʝ�6��ٟ�|&�>��1� �b��j����0��\���f��'�C*՞���,���'��#�H���/Z[s�v�=� ?dw�:���6�S	�nd��5%>,ՁΆ�J����G�����YO���8�ZbB��d��.]��QN'{gD�m���	�2�r@�D�+c;�J����x,��2���|rJ@�� `YOT� �o�2�&cR�w��BT�[�βz-����Z��`f�ĉ�8%�1c�;3��z���%�g�k6��F�~|�h�Ҕ&�4ǞN���|�7�s��-����?���w����Y���Й�I��,g���桲@c�:88 ��X�Я���?��c �qܗ�d���޵�W�̄W@ L5$�~�2'Ǧ��f2+�
����]*Ы�<��$Y�;Ѕ��,�*�**��� ``�A���������~�wha���{/���~�mݓ0O���b����T��,8�Z�y����M��F�J��6��8��Y�| ��'W�.p#�P���� ��8�W���c��
���%6�l�N�����z?7_S���HlJؠ�8-���3li�+D0�'5��3K_@�V�*���z��gӶ<�C�/�pjJ�ʛ�D�U�*�OJ� ������>M;�:�.z[��֦��v���b�= 8����w0���FF�~	���:�o�"�{S�^��Xezݙo��$�)0����܈�h��W���>���f�x�T��
ֵ$�&��ѓ'OB������Y��5���n:��y[6H� LD�b����_eA�j�zw�N��&����TTT�S)�A��_���<` ��y���0�rz�7O��4�,֧�8���f��{��J�-�?�2��:R�7�̫��u�����~f!�3.z�E�v��20�i"*}������ Zi'i=^Ì`��ۡ�*�y. f'<��B������>k@����J�.Jd�(����lÊ�ߛ�������>@<��g]0s�����[]]`�];.����Tc����y��*��B���]�(�U�D6�qI��j�%��B��w{���л�@h�t'~l����+:)�8ۓGLF��wx�H�`t��%�ĤC��Bo���g���ѻ�d��vI���<��B�de[��32�����Z]Z{�z�!��ov��/L�X�s-��{�'E��������fyӎ[}���������2Ӎ+ێx'"(H���T���^�u��.�IzW���1jkM%R�Cw��X�oi}0wV��Ӳ�;���eid||Sq��	Oqo~9���k��ޖ��?߲��%�|Nlz��:���&mb@r�tp�%�����]t�̜&��!;=LrZ�e564�0C�x��t�C���w�`�K=��W9�_�&��i�1�;W��N>���*��#���86,���@4�2���|;&��4-�**��T��g�k�HN�H%���Ͱ#���C�|�'Kh FOenqV72�!���cr�����y7Y����,�ł�%N�)��s�*��]���U��s�i��7/��h=��U�$��+ը�$v �I�d�um�ީ�ק�0�~�3���S^Ϯ�l�eZbG+��˵L��Z�wU�!�[P���	�;�C4g����|CF���44�w��A�o=/ۏ޽t��'�wB�@�����Z���R�E"���buWН��%��=w��GReYǳ���&ZO��U�Ӱ/���R�G�� (�M����,�h����e��Id�KI���ϟ�2�D;��������8&�n�%�U�~m�;�i��e�箻��IHԛ��Î��0�=�ĕK���f⫀�u+o��Qٟ?�C�}:\�+l;x��3����O�����t��$vRn�*�N��贒��u�諠:����땩��9�y�%�w"��|�✓ghV4Bf�Om�-��+��m%6%�<y�w���B�zgaB���&�l��ڬ�4�3�(��m�0˜a����� ZvR�����h���Ԍ����`D�LH^2w���Wv	�N�z���s"������maI�j�~p��K*��y�R���K�x��=����k�i{,{�y�t�Qז7�Ӳ*�۔�������Մ>e��S̭к>.T�:z��cr7Ȯ�8v�A�0S+������z���}ZЌ�d�&������)�z���K,h���V����=�ǯ0RF��@E�v9�S� '���#cc�N���?�@�jU&�ge$����XM��B;1�x
����F�` S
�d�������У<2!�x�6�ٲ�jހ�0���uAo��?��d��p��a�?�hHUM1"�wLj/��������<���n\ȓ(3�ԓ*w��⬮��m�ȳ�=T!Ǳō��j^l�뙟��Epx��Ę�D���`n�:&�
�g�S��ZxJٚq����`�r�GM�VCB�f8d7�0���+�P��ۣ2�l����L��d:��QU�a0�N��Ī`�;�T��<�kW�0�l�3�7��{'|٪�����)��<�o6P���s�v`W_�	��1)���X�Ģ��7������J\�}�F��er���r1�-�G����8�<vQ���V�5@'���2z�RO�L\�s��@O��Er&u�2�ޣ����RO4�r ���ׅ��ݼ׀D�-���פ�M��8��ʙTگ2�-"q4U�؉��->?�HC	��]���;F4v��럍�Ր�
�3� �yx��h܈�&s�X$��+��?�����Up.s� -� �C7�50?�[��M��� #H�o��s�,gd�2� H�BV3M7����b'F��Z7П"��F���E�<?_S#��M��Ĭ��L�D&@d�+c ���tͰ�/��*� ��͋��)5Jݷ�����ˉs�/�rfh8�s�ıQG�Jjev��iZ.���\\���=��<:����$C�_om1(<vkԵ�nzX�tb���2!��٘`Z�ߤ�&��"��	�{*W>�C���"/[8Yv�΄W�u�q�קUT9eBt�N表a>[��j���&$�ͯ��L�z�/¬Y,�R-�p)�ۂ�mʽ0�]�)R�"�����w�Jm����vy�������M��u�j�F���L���0�\�62bdae5vsMNNfd4�!��P�Uo>W�f;J
h=D]�>����+|���0��;:���:>����af��}��ݲadK�
Z	4u����:W?�أZ���%�&J������Sh�RQ��J��V��1b M$��o}(�O���D�?�Td����"1����f)�^1�B�*���x ��̵w�l��zL�/%<�B�\J��I"��io%�/̙�l�	�";��^M�	?�ۆ,ŷ�|C
�dXNl"ͦ�!�_�编s��/�ښMlFcr�m�L-�~I�r#߲s#�~����V&1���0G����IҼt�qR�
(�{�_,3$�?���J���!��sJCN.���8�ķ����1r�u^��m�*J?�WQ��ϟϚG��prr>�*MdAW���U?�V��tU�_kq�ˍlܫ����'uA�����0���M���?�
����P�^�]�n<���K�eέ����Ji~�PK�	q=#CB���a���s���'k��*t���=�zcc��T�[��|UUU�˚1������S@D�*V�e��&���E��u�k_K�J����414���4��t��ݡ� ������ӌ'���^uRi�uy���/����"�L5��Y�2Z7���bB8GG��>#��t~T)UӬ��xx��c��.�'1ܠ�	'�4�dhw�Ǐ�����<�i�UX%��?>1F�/�у�Q:�j��<w��SR�.
�����FƫW�&WW:�X-�������ǩFa�lm�/��$`�9��J�c�6����j'/Ͻ<����ʦW]����gs�,535��k�&{��l���̀��xM��5pĹv�!s��6�ȥ���=π�  @AA��i��5x�3��
�0��J}q���u���L=�g�
	�o�X:����㧄���|��H��>�@��3�o7:�����/�]���#:<�lO\�_S��,K	49L�|'$"(>X�q���@{̈́0��S�w��^^u[��0����O����h��~D
#&��j�W)�	�I̸�`��Rb��-222�EG�(ˏ�ٺC�A�e*�n���m�q�V��:�Ϲ?c_���2��*G<�s��Z���u��~a9�n��`�'?� �~&����s-�%���cgJX .��ci���U�O�ǀ�]�2�<�������_-�z��q������=#�LS7��΢���k�L��Z�w7�^�4L �wEF�u�j�����ELz��L�_-c���g �فzGLP�$�XH�-�	�R0�|�[.g�~�!�pa��ؚ8M��s����Ǣ��d����!���B��[���P
�+�}o�w�Z��QQQ]��]��cG��넳��񰳝l(��n�T���^�m�����*�9���p_�^�˚�b\�s�M�5�/X{:���퓹`4���>2�C��F��OT�bn�a���lԳ���)�а�俱��Γ'OF���
k�p����FD��e���8fMq�@E��aZ���5/�;��,cZ���֭, >3Z=S�OI]��( +
h�(f�(��/�8Tl 3�G��^);p�����ͳܞo8䄈{I �.�@:Cy��-�6�c���q_i���M�{J�����
��'�<[��@<f.��8���6�φVE��l9Eqzn��qs~1�������Vj9Į(n�%��4���r4@F��ss��"�ēkz.�:̾���_GD����v�(̩~C~��n^�f`��W��L��+1R�kߪ:�M��
�p��_��W�d���/��F� �nA�ToѢ�>����l��[//����\9�Ǵ�C�� ��.%z�K�Sӝ�p�?�J��9��N�6�6��F��Lh9Wp�y�e
O�����f�>���l�����$%o��r�UHڰ��߿�X��P�m�^"Ƙ�m5������p����&��+!NSy�+r6����{�սc�a�����"�����t�N����1%�̱c<����W�_� J	u�h.q�	�lS���o�����Jn~�/ej�7���&�eN�F���, ��m.f�p��ۗ3�8���nC'h Zfj��G��v�Y�����'����=���a��pW�׽���K"�`r��'My[Rne0��,�����X���B��qZ�M��ڔDv��=��	�H�Z��p7g'nP\D$�9X�9��!�C9�����E]�Ѽ���n���j�N����AP���l��H0��Zt�(��M?���[b�s�[�8�Z�z�\�3�WƵ��O1v�O2��[C����R��z,�Dq�W�^//QK{��skCj�Xw;[n��?��*��ɶ�|��vG�prd�_�uSu�$䭽A�g�9�g-�͓�t�=��;~k�,N@;��8n�8��N�M�Ra2������IJ<��ȾbA�����  8�N���b�E��~�F��v�0��Q"��Bk=T("	��_�>H� }��݁B������@�g2��0��(a��c���|���+��ߘ�v��tuT������ּt�E;�.� ��w0
��z�4�Du۽��e��\��� �"���,YVY��^+��$&to�ILꯗ�%�t����vG@S�\��_�}�.wwq��ͬ.�ż�9�3�9"�s�e�L(3��֛=�N������q1J��0@;?��+���-\�C�DQ�ݥ��:�xh� ��h�E��
�+�����ʉ�>�2�f��"��P@�酲��7��-��c���?����ܻ��?�y�ϼ���Î4g���KD1���]��o��uw��� n�OC@���9�rjr=:���3v�)jP/S�N1=��DO�#��W!N���kV����+a��b���w�Eo)�j�����#��B�3������{��,�����l��#�$4�A�
|)zr 7a#L.�U��W'~�bS��y���S6�gS��0ܹ��hl[���W�bZ�������Dsg������Ho���:�`o@��z�%yYW�Pl��ֻ��D699Q����.�WA`�sj�<d�} ����B+)*�j�3� ��i�� X�ej������ϟ�8{P�h2��ӧ�D�UUG
��k�V�q%��t��d�����@��Ϸ�i��H�{@���u�)~���׀>�Ud%.iCf/�D�_���� ʢE���3�y�7��!ڤp��y0�~ �ͯ�$����{�:��J��-�'��7�q�A	���v�^�������]:v�I�<�徫:��:>d�;�4�h�� ���;2'ɴ�O�~ �e8��?:�Sy|�����	�_&��VV�LШp)b�,�ߏ���i��@`o���qz��4� ] ?#�,��l��
6�X���G�D��R|{w�R�C:��׮����w\ ܁����ֳ+T��;�� L2s� X�f^I��0)04�8�?]�/^
�6	��~{�
�q�������&�>���$�O5�E]��!\��8ا�=z����<_Z�ey[%�Xq�}YW'��8̠J�z�J�*�/�z�2{�y�cW�����c�m���=���x�U<�"��3ʄȻ������_[�2��X���2JN��/ԋ`������R�`�W��b��X��U*\W���)�s{%�%���O޵D��K	p�Gā��h�wj��������h�̐����7-�Sv �ݓ�fP�lj2ӊ7�1�Dk *ꃉ�o��fy.*��)3 ����𖁆Îl�h�yY[Qq�g�˛Q�⼼o��ӟ�1/聚�95+�����M˜��T�{�>���/�Ҿ����� 	� S)/�.Ɵ5,Cߗֿ�����oa(#	T.�4��ud�����O����pо~�����O�<S�<�~�u��!���47R��eؓ��z�������$��%������E���d�2�:��ս�o��SRR�x�lD���~��unJ?�j�;V�&�g[d`��Roh�!��f#��j�? F���E�>��g��N˻~���)b�Ɔ�;[��Ӄ��_�%u��n"��'6��H_Pb.3��hY�m���6Ϛ�DKI�2= �e����c���_N����S�D릜�mQ���A�i����K���M�>h�<���S�3oW'$�-�}�9�ϱ�	w�{a�R�e�|�] ���H�}=W$_�~��2��'�U?b;�L�4�ID&�E2�9���⭛E��קi�%��Ǔ0q<*y1�����|V�y��~ˮ�ﴥ�Fv���x!�
V�X
�쀇o��tL�yl��;�؈9/��X����HԢ+�:Q
 ���!���Ͷ���|��#��\, ��h����Sn������&Os*Q�:��i�]�o��5A��yÕ��o2��/�R��Vi�s�q=��	�7���[��D�y�i<�@\F�����=8��\& ą`�hF�8�1E�R�2u<C+/m�X��K�����	�nY��l�5[`v�8��Z�G��0V���t��MԜ��_d�N(�:�Kh�?��'~�0^{;��������s����mÜ <�
��̰�'|��iU[4�oI�}����M�-�YK}�@Z!=�Sx4�m�v���ٸr��r05�>ѭg�
�O������E0ЊZ�}�B���U�k�8�㹑F#l����π^�"�egr�"�l�	hY��6�!�wn��yc!ŏʩ�^�����@$p#n��0���O��[��=X�([� ���ǕR�m!���J�6<D��Y�Z���`f�R��td�9�p��	r�>dl�q�8��������n�V����}Q�AKK���!j��kj���٥mx�޾kQ�+�_}�I���XI]��N�#�gNsU*eF����FiC��u��£��jr�Q�+lǈ���E��h�"�WMAp���@�amb�z,�.�O?<KCgh����	�d�1g]�vm<Pb���Ṋ<���(Nη�^*CM���X$������޷��###�a>G�\z?O�)3�AgUx������- �N�#y4���3��8����p[�52���/ý���H�j�nɢ�\b�<�G"�\�9WF�*c��Y�ѩ��ʃ��b�zڦ���������jÉ��w������/�ȫб���Z�I�up#��_C<�u�����Ҵ�z��6k�低Ӭ!U���廱�~q�����z�Oc�ŗ�m���(���0�N�� 3񀁧���}�ŵ�R�)V�y�&-L�m8�i������$*&& ;;�ŰO����R@}�]w��İ�N
�n��]�cw�d,Wl��5�v��s�+�?N��������)�Ua^���{�� %��ςx`�W�ZM��}HTԏ��\3Pr[O���S���U11�0Y�nl+?�/�@x,y���-� ߨ��鰩jN���'������eǭ�g+KO�
7PR���n�����J�g-���Q�45��6˱��t��Wa���RϞ#ܟ��������>UX�gEv�W� X�:aH��a���`	~c">x`=p�g�&�ڞ> �	�:�-��A�\��Na����S՟=vsF�<[�-,:=��6A%�az���Gc2����&<'<�ޮ��_{߲W,�&���շ����|4���*�cy���t#�f�g��/�x�8�z���_���� �'�###?�-��Y���l�jP;=�*�v<�̓}oA'�
���@ᕣ��$,�VGR%� ���s�����a��5��0��>�q��5�7�M@p�D�~Q_�cTXZ�l5<`X�Z]Q����Qv�a�wx^g�?�qg��b�+s�A-`hE�z����j@d�����j@񫘣���]E�wov��Y3�Ȏ����XJ3�U�>O��;W����f{��uZ-��x�bn��s�z(u[�n���^hom��̶HBMd����J�ho/�m%�}vp*N+�*44�p��>����\���F�egV �5���c �v��U����앬yQ�{܄�-����M���9d������P�òFgi>4�\���������B�a浄�[SG��jH��k�\�3�=����>:~�ؿ�g_x��ׇt\M�{ژ�I��7(�IQ܉S�X�m��p�.���ھBEM=�I?3��m���;F�)���q="�~�ds~(OB7��~O����@�Lu�����XZ���w����*�T���`[x������g��n���:9 d�6�3Pj�'}��R;<g�KXhH�_�pE>�HT��/��Y�1
�����Ij�؋��5A,VP��Àv"�g��Z��B�7����>��tv����I��5)]����hZD��	�^����[�j��%o0u0�䩿���v�N�+�?.��?�xý7P�\�%�ݳ�)W]�D��>��I�*�miQyg"�˕�J�B���N�t��UfN�gI�$�5 D��p�K0����ik��f��l����nG�eq�1�-��)-3�i�q%�..ش��׽*�fS��k*+%j۞�NO[d�Pd��$�
���.�MU��)�5]A�j����9���}��h�1�=�k�}˘Bm$�W&��Y��4�%n������Ş��v	���{��m����}=�}��b`��g<H�e@�[�JU�M\)q�Tv�s�N;�k"{J��>d��v��vw�qY���*a��v�;Vwm������Hk�1�5����z��&������Sy�;%zK�(�f�~�遣w��y,6�����وT�줹g;J��R����'6?x�^1%w,%�쑡῵�����>�.K��K�Y��`�g��[��:�#V�Iɕ��'�\�8����466���-�����ǖ5r^,�,�����b���K=t5g�j���E��`~c�	��}\\��O�� ��>����1����m�.�ˉ�����6�1V�%�����PP�V&,Y�()	� ���@r�Ֆ55�=p}����$ҥ��>ǧQ=rZh.�����	�lѾ�	8�d�+g�����O^^������!9ᐨ�ҥ�똂�����:���������[����WR�dk���tt�)�-���g��T��[�e����c����$~I)^OAl$D!P`$�ұ�Oh��r�%Ay9sO/_��(���ﺪYrr ݛg��M$]��t�:?f�oĻ1�	����+��K�z.x·��t��J�Q9��=�ug��;�H�`��W]�ex,������U@�*ym��x�?qu�Ǖ�m��rk�ߙ���i�Ef<~2�꿸R�`gjε}�fo6� �J���pWl"��ʪ���[`.�����������c]��[��	_�@:�b�8���)�2������}��7���^��(��_�ԉUN?��ݍ].���o9�����,u+��5��8���ֳ�6�͎O�y%Z}���]S���H�^�����n�ߛ#��ʔ���p?�8�_�X����]��8w��JJ'�H<���bѼ������\�%N�X��. �>>9�E�T'���\���ԍ������U��lZ^����Pq��$�/�_�F������͟��ܹ<pb5Fi�.�7jV�j0��\$/bRp��ĝ)\M����Ϋ&K����@� ku���>jqā���.�NCj�:����f�ڣ��wK	�����+)���w�b�4t=�|�|	C�z�#�m���w���=� ������T1\��B�{��T"��	/0���Jb$z��������]D=�����ew�0�O��!�p���/<W�=L������0�+�,���/���=j?;�ů�NcCÛ�3���NN � ů���4}�ۏ�����<'7wr��{"_׵LK�M���Kx����}:���R"l7,�����'�m�*�.ۚ���7wM��N�}�����Y��`Gg��ҁO����|��m���9�_=r����o7\�;�,JM!��-��� �b��=b�(vd�c�]8��и+vĀ����E��m�� a�4��K�i����W��k��� ݾ=ؘ/��s;IzDb�OM�R���>#'W7�q`�o	 n�z�������f����e|{<��N���{������;������8E=|�U߃�\�m�6N�$��TU�}�h,��n�-^��9����c��}}�����v��Ս��ȑ�!�& ��^_��Ғ#5�lW!�5n�T㹘=Ak����m!ͱ��������
�~��= ��[����y�`��|7�zc]I��3?���������k�ց���u�,�O�����B�b��J�+k��W�����}u{_Չ`�ǹ��9��s=C0�r2�.8*�P����O�w��O����z���*s� 50����H]�<�Y/�o����_|k�ؚVŃ)��J�.�M�瑉i��`0����`��x3TC�.8ܪ�c趙.�b9t�м?��l��jC[��}�CQsppLH�t�y�����Ħ_�x
υr�	֑�D��vR��_:�9����~*x��W��*+˯����g��f��>פּ��'���͆'�k��:�{Q�*%���U==ZYY՛� ��lS>C�櫷\����i��o���ڵ
�����
�K�w�����k��K����!;?�
��T���'+��V�[
�xܷ���-���HƵ��|ll�@��H`�H�O*��z���}�ug��V��D���uuu	���*M�O��r����M����ƪ�����ش35��1VG����d�f�B8�[}�~�F-Q�%��FwNCG3�*l��o�f��T����������*2ɍ;���<	��6��=Pҹ�s���Ͽ�/�xɞ�k����}{���Tz��U��*����62���eQ@+��Tھ�W����i�	B)��Fϣ�yt�bLɍ��eɸ	e�;ӿw޴m?dZk�̄ĀVC+�R��둂�0��PY�p�Nccc&AAA��4'@iR�|�aW�㱐%�n�9�ԅ�?��jFB�9��jd�̤ȝU��]lKMr��pX\�uX��53*��:z�<�1�k�I��"T���/�5��+�����#��Qe\j��G�u�S����RJE��(��M%3��)$[��TB6Gvv��8V�N'��8��>2Y�������;��^�^�����w~>����Ox#�����st|��ق�"9n;w�g����{s�=�q$gW:�N.o �q�GJ�_��Rg��<��t��S�x���*B��׾���M-J�K6�o���=����u����q��U�Z���h��u�M���h���2�j���J�vފ$�R���Pq���  �66�#˕�#lD��=��m�%��"�frQJ��x{�l�eE��c����;/�t)���4��r\�{�"n��D��`5�(��wWfo^(%���ѕN�MQ��+�g���YYY���e��a��OMC�������[����&�������K�h����^I�+����OVS=ބ�_Fߤh�	A���ܠ������+C���I�t	��#�0v����M�=���bEA^�^��?>�M��O��q��f@�L�&p�.<�x�M���gV9�j���Z�_�	L	��uH�.v�����^���~����Ǽݺ�J��Ȟ���8��~k�-�Uq`z���˅Zy-KK6��G�\����XM2�<�Zyc��K���n�ߩ�;99����%��ݪUSwp�C��}(D`FQMt��؃�&'���Ϸ q�W�V#��jܻlwoOj�6�	�"0�VǑ"Vp�s�Ǿ��F!�Q���;Q�� �����E�6T���E?Ju�(U�fXŷy������l���}�S�8�ھ��+�ۛ^�!�H5$�lR�/�"��<�/^�p��s#��(�<^p����77��m�۴�]��y����e�Sn��{�a-t� �3�{�����#�}i�.�xЃX7���[�Y	��:xe\Dcs��(Ɯg���&l�Y���{�{}U-��&�������T̹=O��P�^�5h#��}?`�������#��n���nC�������c�����K?wZ���\w�m�:��<��
��p+\9�~�ɀ��ɾ>s����g�{*���o�á��C.�/��&��_PF�D^
e����UI*{鮛��uW��~Xhl�wj����u�Z�B��Ab��aW����R�*$��.\]}�t��;�q>>r���֎Z��s�f�?y��2뾽����זֵ�!IJLE�yP�:�ء�\{��R�*�7 �����MHP�0տ�������x�'�1ٗg�<�3uԖ���6�Y�?ˠ���ɻ��'�Bw/��6���v_��Ʉh�;T���W ���)$D	�ܓ����@��cd/��)�з�`�������Ej��SN:�W�l�ΐm6`�p����q_�MZ�����.OwY���Ð"ᕮ���'.4p�K6�-L�e,�~�5]����9"$ ��C�5��b{p�,0tL�E�[.B���oH�С,���VV׏�Ԅ�cM�?�U�������=?�w0K�ų�m?��p��6�� �$�CӬ���4���\�#�z���ԺI�?�}ܪ�ېF��}���<&��C1y�ϽA��V��T���O^��@�)75�*���+�"%p��	��/���虼0�+�'�k�(
�*�~�%(�o��ж�Ѻ��h�'�Ȳ��hr?�+Y�y��ၰ�\��1��0��������`K}�҂	d�|��!�)C7C��6J���g�C�ʙ�����˵ �����x/�ؿs,M�X6<�.R�O���$/a��Q]��<��}�as��µ&�HHZe��EM���2;�.��U:�zFֲ�߬�Q{Dz~����݋k��p�Zԉj���Qu�А �|��7�Q�n->�%�j�ͯ������Z��S��������!�����������Hf�ɡ��
��rB���QH	�TF٬��K�6��D{M�_�'a�9�y���e��9X�̎��
�^�+��X���:= $��$'��vo�^�z3���\���ׯAjI=�BcD4����?�X[7�g��:�M�y,޵n�E;'�X���f�pOY��z1���lF��q�Ĥ��G��KJ�z��]��y>�z*���7u A��FQzq�s� �Ǔ&�i*$�)ڌHC�]\�sc�'Ap������D�Λڐ̒lH���͛�%&�����V0����j�ޅ��>��'�Uҹ�
���$��J����A�R�.��5 ����O����^m����??��6X�~1�+�0ul�ʢ���`bZ.���^`�L��]�RN�cy0�q��2	��R��Mi)��� ���U���Ь����>��-4N�5��F���8y������D�L�$i����e�d���5�ى����7���Ŀ�=!�I���=E����W4��ʨ��H�����⍯���Y*#�z.+I�>�߁K����N|���Y��X܄�\��#������n���i.S�|%֥���7d�f3���ms7�K�~�c�����osA%��ٰ%E�P& 7h7X��+#Z^a����e�<�����~dM?����5��r=����BV�D�߁M,�+Xӟ��!/+
-%iIl�ȳ�S���29�O�W������˚x�>�L "" ��a���D`��q�x��l0'�r����:IL�rS�2���>W�� 
��3ȶV�S=���C���P�l�ϻ)c:�R��P���������b<�S<o� �
�� �'������2�Yvߥ���2Jm>x�����$��)�3N��T�;`�˦�	 ���.�;�OBsR�Y�/\��.��UGu�s�`S�vE���,2�?b(۟ˈ��ʢ=?����K9��:P���)&7�$�oJ�T��[� �yzz��ᘹ ;��C���d��R*FF.����p+���Կ�tz�x�`��|�� �o�Ѕfs�p�T�޺ ���i�����\bp�V����K��ڎ�o�y��ҳ#��������0.R�?~�a�����ɤ���>��O�dR�[����Ʈ!��.5+�_�|�	�*q��]����?^;~�.jL�6/������U��Ⴂ�囷���1�P:�57
�ef��Z�Lp�����N�o��1-�Dq%��ln���Pd�S��ı~���7y`�,T�_��n�,�*מ��-:n��%iS����z|+ 	��1��_���gil(6���7�.�k� ��T���o\��Y���q�l�rp�*Ɇ
S�H�JuF[�ϼdl��*�n�] ��a�.B�8�[=
I��V��*�Ĕ�e�}}���@���,
�!�W�@ZF&f�+u��BɃӣ�>��U^8���ZN��̆���
�����k#��ɕ8]�����6:�˨�N�о^,j�$��쵵�>�LLP�2%�-՛::�}:Rn��-�^ݟ0c�X�L� �]7󳃰�'�X�����$��#� �kTa���@��掱��g�գ3\���0)�����j��TU
.y�K��Mz�h8�����tX8gW�5ԣ�V�h��V��e�{�~(��lt�e���y>kzGl�L���������,U �tf�f�����&�� Uo&8.83r<M��`6^.��n{,�iO��a_C#�B���U��ك���߮߭�>��(����5~P�������\����_�Y�
`�3H�ٸ=��"ָ.�:X��2�;�L��/�!�����|�ϼ\\m���lU�N�oũ��{h|�i<^�u|a�7ċ�zmkۏd&�{����ڏ��7����6�bc�a ޯ���p�W�ߪ�$]s�ĥ�A���C���nt�2O-n�kj�kE�8��L;�Ⱦ�|]c�1�c�]{��۪t_OO�l����q}|�M���G	���*º�5cIFI�D/6nY7�=[U�;<��"��}�!�8��^2�g� /ǞM�~�=A��Zo�׈�J�9\��TV:�<��j�+��i:4�4�>�r��8�.�*�0�d��u7e?}.��B����qG���l����ɖ��;ގZN����2Ӎǃ'�	��5�b�ԑ���s_�O��m��[X$
��I݉n|�NY�D"�h�~�����Ǎ�@��O~��7��]�����2z}�>S���Zك����]���[�(�������A��
��Ƙzz�bkfS�Gg%�����-?�F����	�@�:�=��*�������<Xo����\D����4J�5�o)� �6X��t���\���-$}�סNZ��Ĵ�ѣG�+�1�T�srS�?���/\��6?XS����3��uUA4E���ۆ0��澖ϼt���h�.�\Sk�
�=:��)z��6�ֻCm�P��LJ�f8Vp������:ɡ�M��M]����c<�Ht�|��P)�3Î���>�q7��c�\��y`Ԛ�T�.�t��=���ω��V��x|q~R��c,R��,?I��vee��Azl<ӎu�J�Q�_�(DX~�y,�h�>EG-f��C]�cЙiЧ~պ=�L�Pxl�����@N"�ߴ��{���TY���%�"ή�/�}�}!����"���\�>xn�B�SRP@g�7L��A�:�r�|[i<^�����Y�<��ή�hVj��Ɇ����s����s����6X��"��˂���Z G1FA���A_�m,�={�U�j�}v��r7�qo{��m�+T%��W��ؙ_�߆���e�=�*><;�g�u��b������,2�˺ꆻ=�q:�����8J��xe�x��D#�W,LF"0�K`�]�+tR����������?�L�b�g̳�]��_�F���
Y9��9z�в��.Þ힄���6����Y��.)O�xg��;`>d��&..+���ee��8\\��ν+�ԟ����27�Z�<���ZZ��]�3�w3q"�)���	$���3x{��Dئ��m�T�v�����KLBL�]n:o݀���o�h��ң���ߖ]M}|ꋎ&�wl*�.���,���}��:������h�S�ǥ4����R{�!]Z�&�ΐ._E���&�!�y"��	[\�q�)�pCx�����A��Q6�Q,�`�.W�����B����J>��^�{}*�|������
l�ΓC]���T]�;L-�Cd�D��B��\
Ŭ��cR�e�;m��]�S%\O��8���N��+��oۀ���=�S����YiI�Eǖ]��D��/���QV6�Q2���Q{S��^FF)���{oJ��E8t��C�2��Rgq�w��OZ�7��i�� 0/0�����הL����6�j�U{��'��w������(^D7�{���%��1��'��m=�ZMPL��C뜫F`���V��ޯ-�v�`��8:m����J{,d3��P����c�J�p��.����k6�U�_���ݗT9���y~�B ^�C�+��zx��2���t��2N�4I��r�6�|��ڹ�������V�<Pι�QNy�N�e��@Z�yF��,����mt�)0	6���f8��	���p}��v�#��d7��J��+����#]�(���{����˭�$!4'F��wm�"_~tSi�'$_���}���C'w�ax���ϥ�C�����y�~��!��������~]�H^�6�����`[W��O�ݫж�l�����`\*Z�+�DÙ��M~i��2Sv��)3�����<�g�?w:�s��ﷰ�� 'K�)$��.�7�z��
�G�g����i�u���G�LZĞw��mx�������j�����F���.U�N���*&c�������j�Mt�33A�+(��'n�NSS�Z�4���ף��Y1����W�V����g��BZ�R�*�S��̘��MFL�Bb���ɬ�[�A����:�M�_`�0��з,���<���nblo�\���?g����˗k�4�svn�ݙoiwj��C_����n����WPP�3Z��;����lM��DvA|��	�x���P�w��8�ܚ�d��4��j�L�Aal8��;i+kk���k��ƀ]q�<�p�z��9~nQ
Ӛ]^^�.�R׼	��}�	���2WCK�s{�����!��b�LU����܍��)4���]d�ѡP㾚~�\����!5�Y9�0���R�}X�щQ�$�\tG/V����\y�b�n��/$�����*���(e[T5:j`ii���a
L���#B���@ 0{�=�Ç�>�4

�033�s��?���`�c���I����-���|���>bf����
�8,E�W彼XA��J�ttt��ř55�'҄��^�N�����H)�@�( 8��A�������O��`K��K~4�ֻJޖ�L�{ssӒ!��%/&.nю�澾>��Ztqf~�=`w�U�4���-ml�1�XTr�GFF����R�l^8l�l��t�s����dc�T�,m�6x Hb�$���40�~���Q��p.�E�[_o�������t�y2�6���A^_?:��q���"R�@�]Ee���8|�s@k���gΜ�,,Tq��|biy�
]�8��,%e����R�0�ǏǅU�q�.U&!���r�=�Z�V��זʐ� �`���f���y
Vbs�w4[����=_��{D�5�n��eddܡ�⾛�lkk�Y�Afy����8�׎��No\��]�
�-���ǘ��+ٶij/ɹ ���#�,3}.F.��I}x�wl�qNy�B��N���T|�^'��{{z�'��Gk�댊���'���M�ֆ����?�6���� ��w��N��qQf�S�y@^gΞ����U�����j=PW��D�kj�bQn�VVV��W�$r�\��#��U��M���� �u�1_H���Q�u�,���r���6�)��������V��x��첲�����}ǟ�0���%�	B �7��㕿SR~��"��X��t`�8�k�@�����U�CCC�1�S.m{K�`�/:�0nK^B��؁Ϛ���)(�0���ٖz�� t��8�B��7�J8Y��ںChĞ҃��~��w��p�]7�fn<��qs�\���o�?���yu�+U���y��M����_}4O{�}2PC;��=�}O)�7W�'� ���PTD���A��]c��Q\9��H���}#e��¶'�+A�|u�3�!�fg��.R���E���{��bAu��������� �2��U$MANE�����jZZ�=��� �k}�0 �
�i�Լ֣rOD�0[e�30��x��?2r�;N	ܻ�A��+��Q�?n/O��v�ݡ�CU�.$2��/O�-{���Q���.X���d��!@%����5Y̥
����hM��?Y،�or�i�l[�.!�dC�\Hs$��-I`yUբs�ξ�S�2S�����	������+�0�̫`�7��������}�>���-����7�b�e~���]W'�(�!~��%5cc���
5��`� L��}E�� �*j���v���eA�'''�nl�g8���>?±�ۘ$������
��]S]�h�WL,q	v�]V�]���h�&���Hxm��^
o���UW���PY)h���cr2=J����|gG=|�����<�*�Ȟ�z��p�_#0V�;m-SO����T�W��fF*���s]� я��ǰ����R��h~y!r6zdD����%�k#�U��Ouut�Kbg����;w� 1���)+7WAi@��4Zq�����72A ��f��e��쀮����06�LO���	��ny���0^�U�G����ʿTU��Ӿb����{� l3��f��6�5��	}�]Uj��`�Ż�����q��/�����ۺ��.^A��~e0��>��������w��L P�j2#��PM��H�� ˄:=1]TQ�i����w\�V��E�,�r`�Ƹ�T�"t8�˹��˝fU����r�C�	�(�摏�IL��+�~��]&S���q�h&��$�؈�>x뻑�����5K�jr����lr��Ν; �M/䕺,jem�PS�]����yo��UyS��H�}y�S� �똞�,%z˱���Y\|����nA �e K�Z��Pl�-=1��hhfFk���߾�P�㞷3m�%iˡh���~�6%}��������uϒl������ɂ|*�PB�\�����aj���{�0Z����U��; \��M�?����,�'�5���ђH��SƼ��cN��b3(D|g���Ǎk�	%VTU�����H,���K<9���ۖ�R[���YJ��#�C[f��b��?�}#|��9�Mxx � ��E�U��\�_%�~*9ۇ䂾�	�9�Z}��9ܓ�A8JG;o��[��C�4���3�I�����w� @�Z����C��B_Z+K�sj1�"����Y�@���	$�r�*uqu��fk�W�r)���XPU�k�K����"V$$�	_�?ت2�W��y�V<�����?�޽{��45Y�+m"��-�\�ِ���=~,����i�Ե����0�#��Ƅ���_eW_��OT6��ݱ='�L�������n-V*��!AG�I�&��5��U�O� �B'D���G���aX�$|�fm���������0g@@@��O�z�F��e>\�>Q���6��+ �2u��󞘘�}��l`�k��M3�
JJ!𑮮�Ԅ$_�	C��+~���@g~�8�.��:��&��Ę}��@�v�l��	��)R����=���^?�WSSK�:  g�^�=]C �K����s7XϹd��ɰ���I�.N..�N7��7n0~w؆/����~�^^�I�=y"�{���B-Vr+�?'�0�|K%ءH<���b/=[��T�A7��z��������zXsY�J6t8�+v47�U����s0�{��+9 cǠ�Y�ǡ��䯖.l
޼y��1U���dr^�\�tl? ��U�'$$ĠN�����(�eɶ�Zn�]�,������P�s�]j �(;��aj�Ŭd!X����>o�=�!zk���l��	����1�hLt�₾��[ �U.0�D*��/a��Q]���b���ѳ2F�*���i����r`��d�M�KJ��D\:&��e�)؊�S'R��0�f@�t�z�
����r߿��i�jت(�P��1��[����"�G%o?�����4�p��M�W>>>֯ƣ,&��]\\,�/�
��{z�Ԥ'.-?y��=@*�M�EB���O1��-<�,�`�svqwtV�mwk�Ӛ#LK��U��aX�&�|RZ
"���\Hhd8������C9�C@'��nB��Kͻ(�*�B� }��a0��Ȯ�(8��i��$	/WLx���x�k�}


3�{��{{޶��i����m&�i`�P�!�Zsps�-R}��h�GJ�C�=���9Nr���UE:�L��%}�s�#)�>����D� Y��+���"S�LnTcے��T����O:� 3r��Ŷ�\�I�������5�Yo�_;J`��u����&&�wk.#\�Ν �/�=~A51����Y��SSSS^>��w����J�����Yv�F������$%����Έ�j�X"쵢DKg�C퓯��צ�$3?~(�[���	ܼ�V᫢6�g[r�Q[�z���7ɫ)Xq�(,?ː��K��<e�}��KY9��EW36_�n���n`�h~����9Uޱ�L��ɇ�z@c˕#�++q�ui�-��un�J�a&�������YJq�%��<�Y�v�Ω��&���b�S�l�[}�%��9� tb�D%��Zu���ZὙg|)�Y�;�Ҡ��Gi<N��q=/m�C�^�j���%o1��h��av�ª2�U�H{�'a�������0u���h�\_ggg9`4�´c?'̾U��s�	拻����2���L��X�s=O4�>����X��54ڟ����h$I�EQ%I�
33se`Q�ϗ<C���#���`jJ���p�\	rrr��m W�u�>��sB`z��3��XG|@���||�SSS``W
KO\ aHHLNsB%G]O_��?�m��N�v��5kna�W�������b�qϿ/J2귘^�p���vR�
����ޙ��!0v4���w�m�Д��3YqFQr�c���>(BߨG?� �p*��g�V&��0��Z�H[���}�B ^�ms�]]\��S����	�=�7D�Z���)^l�2HN���O��!�MLH�*1�\z~��)���*j��B[�-o�'$iX���)h�|W���wYS|����#N1x�;6x��*:ԃ>G�j�!)(�z��<���Nj��X3��{3� h:�fv�3@o�����ڲ��fX��౅E���_ �e��x`�E%&�ْ<.�*)��p[n]�B�f��實���'%�Z��ky;���S����.�j�O��
\t��[���eg�:2�n R�v�@���up�Z��㮑���]�2�+-�3ч������V�q���w��sj1���O<�����������KK�jB��11����#@M��?�T����*1|�������ʈPx3������r�I����,љO8
��;V�ŕ�L�}���������L�1$;�r���^*Bu��%BG��o1�d�˧.IHH8��゛�\��<�[�*�:�s�f
�[1P�X�����1�T˼��h ��F��lkkk� �ް�~`�����[ECTT�Z 4� ��c���!w�0m��+���Gt�C#e�,��
�Ա��S�w/MzM��&;����5�xIsR VA�^�y��w͐5߰�a�JI{��0H��r��D��5��y�+
��3
�w0�G�M��ﻮ�����׭�~zX@�aDa!�R��d�g��\�A��{|��ѕ�}Bbu]]�.;�D�U�v���eb��ŀv�b9�����|�U�y��KL���rM��ҕ1�<��Q������ c�"���P�3R�����l$E�����!����}Vk�o����2����� �	�͙3g��@p��ac��^.$0�Oߋ�����Wϟn���S�'g��m�h�KU�8*p]��B�����e~$��+���1�v��6�T�^����z�~�U���d�����e��-�Ȃd��^a�T�G�	�u�����U:��$�S�S�����f�� �zx� ����A䶷$ �j���N����Z�!|�΁<m�7E�+W�J���*��#ߦ�2������Ѯ���V���p"t����h���
��P�L�3�0C���E8TQ(#/e�zJ�444D��O1�ʜ��|�E4N�ޕq]���C�ll�������AZb�8v�z\�ɩ�������<-�_P�n���U,E�lL'���Kt�X#TPX[s���ͥ_�9�bQSSSu�
�'%ţ���+!��|_XL,q�D�h�7 55~�p�Y����3�!G�a���yN�2��͐uQ�c�t N�R�]W #JKKi���^ +���;�XIp+>%���딤�kTa֌�O��{k�!�*4��4r��V���|�$"Y�M�{�Q�>pK��f�i�gYYT�onnv��eA7�$؍�׊�/ʎ��v���4KEz�{���qm�#������B�.ͣf�+���j6S�`���dq5��rM�}65=&��8��]йg��� sVVV�>^���RR�@i�]�H�������6�6@� ���Tn'
��HCڥ�
]�Zzz�6�����g>��:�r´��o��\���$L�;8�
Unzk���94�hG$S�_~u��R�Y���B�	��3g�f*DMMm���>����%���ٙ���&X��4��� L�l������`nаj��WD����[:���'h��)  � ��0�=?H�] ɚ!S$J���-�&A�+]㉞��1���zz�LF����ssOd�����N�����aX�)|��Q�R���8ѼM0���p:���߿����*�he�ON��@���e����Yd�QIfay96��c����+������⫝̸�[w��JU��� K��]��0(�����yYZ*�z��FD�ͭj��Z^[;n�֨ԥ�(]�)�'��I-��4:FSl��ƭ[��+* �}�}���(��A���6ff�<������8�l4�5K+�(@�������b�tu��"���fdRu<��q�~{�q���/a���}�@(��|���q��6�x9ɃmS��}�ОE���_#����pj���c� j�s�Cs���!fj
ΖZ����7����F ��4/h���&�Aj����M���1芶�1��]�0����r������r�LP�T�?q�/L{cc1*7�/X�����}�k^�6=P��H�vv���z�ͭ�b+:F_�sEEE�O����=��&<�z��mv]@|�j�[�����	,� ��(�J�o0����m**� �cee�	�6���[�@��l�k�0yfq@����S��E�KҶ6/^�(/'���,,����/��8ඇ�K�Q�"Ҋ'���΢3�lTe���z����	�w�ϏnBEV-�Yu}������lp}��ff2
\�\�_��F���=}��Lןm��f�f*��v��%/k����SՅ���ܹ��eK��}�穧TttІ���x�<���l��Fl�.1))ڵ!������R��]����U�o��S,PNCL8���^�l���BSӒV"C-*�ߝ/q�%�$*&V��4�krM�!"�`K�[2�DmD���4*"1�������2KZ��$��S��R/��Δԁ��t���#/&���6��֑]���ԛ�I�����G;���ε;�!=.�H�0֏�3%%�sE%�Y�KZG~ˡm�v9b4jw�*��k�򼋸�I��xf�ًE�
���C��[p8��5������dn�j�g��n4�ޤ����Ɩѷ�O+ۊ�T�66�|�kn1U�i� ���̆Psbb�f��d!-�����FΪQ��n���&%�ky	(++�}�C�C;�Z����pBJ���?��u�	��9�eqs����ƀ�f�1�h4@[�e����_�<wFPP(+}��b���UY����:��iFG�m�=y���e��>ꞺK7��\`�}�^� G$y�./M�\���9%����a9��_�!�J3ӳJ̾VX�����,�T�o�����	(�
�����Orm�7��F|�@�Y3������Դ�d�E=��ɋ:K�ϼ�\yQN�{gz�V�RM���c﯑;�	Ӯ��C:��<H���cS�،�;�OLH:��kT������co�MW��}��;���O<L�ju�&�@~R��1��/(�E���j�$�p@`�L��y�+�RQS�i�ο�U����G�F�M����j��w�Ѓ�/z���SZ��ؾ�]� 6"P��L�%�-L^���`ұ�����*��˓hdb>��M/�XG
�@��4�g��	g������0 �ޝ�$�Yn�{��QE��:'���]�0k��"��G�3�7���!� %߹�������fC���!|�.1��_4�[FW-ڱ�ۑVW���G2������@E"���q�H��
t>z��y�z�j;� �1��t.@�$�һq�Y��
�X�\�P��ΝE7p�~���V���9p���p$Ͷԓ��R�NI��oP����������j@���~����f��ʙ�4��Н��5N938�x�ݥ�2�+Q�X�=\� O���e����R��������%@�!u�~'���钘�?\�U	h���_��y%��m\�ЩQ��x��w���8��2z�o�pl%����3e�+�c����@��5������i��C��Bf��I�U�M1�w�(C`[О��^���#��� �[��WW��?e����l��A��d!:������Q�[ ��O5�,.�\u��^�2��!��EJJk���)������?�5��옧��J�@8\�N�(E8���Ã}�����/� 	%�-%��VSp���#H��[o���7'���ɪ���õw�����|s���+螺��E�!㯼1U��!�e��Sb�!̻(y&e�0/&!uM �)�g��Ɍ��99rPl�_��u���3/���;�	ͽ��j�xG�&�Up݃�S|||�����@iD	T�	�E�,}��="��W���2�`��� +kk��h����j����$q5H]�x�V�#������9	m���;"%p6�SE����洀SvZ��4���y��mX��yԖ}5�Z���H�;ą�%w_Z6��&º��氎�yɏ�Ǡ��Rgi}��8c��X��ǚL�w�l�������]�	�?��O���ݻ��y���>���ө� `����6�u�����PV��o{	�}�r?�����~�"~���P����AQ���p�b����o�n�V�9@?�@|�L
9��4���0=�1 HCУ��hU����`����T���� �������ڑ5l����~�<Q�N���b�����S,�7�f ~�	�{:�Q	�-eδ�>v���](𨥠,�����HpJ�t��~�����F�ƎN�������ɗ/_�P�"�������$;�+�\�����MRVp�]��|9"(��v�	�hL��)�i 	+f\����4����J�����^
��!l�.6z='��!�/�2��RsXr��Y>���u�(�������ͫed�����XJ"VT�;9�~.Y:+2��V>V�y#�/LSej��������-BK�)J��o�^l�	B�kXX�TJC옗<�rr殮Z
���'yCQ���Hڅw���e2x�0n�5�j6��#w�qs?"aT n� X�h̦op��u��2g=0T~ڢR�j�ͅ�י�^P���^[��_���7�#.>6��!�w�Ssc�f9X�'u=Ch�W�-�F��%�`�i�>k��\��^���b0!�,X���"��G|������3��6�B����Bծ���ܸ��%F�ܼ��zQ�x����'̀� r3p��>�ٹ�}�j��2�y��HB���>�ɘ��h�aȘL��
p�P72��Tx���a__#kR�t��{Ν��(m__���w��i/n_	��X�~��D:�  T��@���bfy9���"����n���W���T����fؤv��/[�ġ����b0�N߯<<q��j Z=P�/�����jt�9�|�9�`�Q������q�@�i���q���7�
s�\u�3����	ܒ��$�ٳgK�u�7���f��Mjy�h���Z�z{�W�c�lP�}ea�WK��-:��(���75ͨĐ>d<86fT��4����c�x���t�#�����*��T&$y��L��l����/��D�d��B
�ۑ�6�
���Ϟ�rkr�m��b�ihk+��?0`�`H����3L����DB/��0]#���"1�jQE��;����Z� �=wj������S��f8j�����2��M�=�B�N�s��yG�8���d��5�)�琭��~O�>�U��p@I����� j?-���-Oqz15dVIII��d�������
%E%%�*�j�#y)��L���WAr�"fps�[0�R�d��Ah;]ۣD ]��Ȝ�Bද^�������;��B5#�C���44�(,�@@�=���p��)��>�[�� ��Kl&>���������ǎ�	�;99���9M�l��������R�E���]�� ����@ ��YY��W/���>d2zhn9'}�0�F�����s).&&F��Z��]��xC>I���[T ��iu~���>�	|��]p�9bt� 2W���q������"۳���J-@���� J}�ޝ1��'��B`� {}�'o��V-��$GL�}����ӣ� �p���	*�����oU��9�z�n�R�PھrZM�*Y$���se���::���J5��B*;"MMM������חڏK�T�����N�����|fer�,>!A�ȍE�m�	���_� <���?u���W�\��,G�4m��.l��[�m]%�mj��H�B� ��6�U��V�S���:��x����.��\h�@�_�H��m`;U~�U/��=�~ku�K!-�^�)Qz��Rmڍ�4Ad,�I�_���^]}�R��OOVMx��dK�#vT����1>+"Y�,��Hr...P�M�Vpi)�5��(�=���1`e[���'����)T{���A͏ ���aյ�XUr���P��)�b��7��!��0E���x\85H�&e_td(�^]�uWv��e����^_LVV���˞�M����[�ku�������&���)�sձ��$}#�q2��nͮ7�oÕ�(�^v�1Dw�P�s6�^���ia�[�������C���ܓ�O������߭odG��y.���4���Y֛�`o�n�)D�S �����wR�ڑ�ua[O��<����]�|ӁR{iP;Pj���D�c�GQ{?0����Ϫ<�~2�T��9%��ڛ�(]�x_��bh[ڜ�g��z��췧�E���QQYy=/�=H_���G`c�<��3����s�}�X�B��f�N��Tt<u�8}=��� �b��� Mkrrqu�b�ff����4.�J��n�|���;; Fk�n\�O4�hU�J��BJ��|�YJn��DeT��V߂��9'��fq��ZdT}������j)��Ը�m��� N���EE�!��2�)à~|����T��ږ�24b�WI�� �O��>(��5���IE��*��n- K5��1�2������f���X���nAZ�����(͟�`	�t��x]�g��v[\���Y���z����-",H��0c=��\���f��o����/��B#�H�|�±���\$P��&�so1ө��������ﾭ�8�?V��G�������gU47?���>�"$�~���eSk��/�E�:#�������Ǎ*��O����/,����.�cw'�������������-�?�Zш}� O�^)ԯ�;����W�k���U�G%o�~���֝��b /q6[sWd˲�yxG,�8u+��i�Ն�"LJگ�|���Vn�JBA��JGR��g|��܃�O��0rg�!�#]_[�Y�!#�����dmnn^�*����,e��,�����������ϑ�XŻ�9���e�`UY)h���P�9�3.�ff�_�;?d;��\�K���B�J��z�,�}���"���tbb�ז����;�Fcw1+�9�c��h�l0���(=�l+�R�6~e��X��{%�����/sx)+��(����"\�'a���ƾ�p_�;�����W���	-�4����8f��Z���Ƹ�����C�~�@���moW�;��sg6ҒN�c���:�s��\�1)���	�Cfc����S05Uh��P���j�Գ�¯<��ا� 4N�����ڔ����w��U�������棶�JT$z��HUe%�>���\�6����%�4e���NB�6�؀�II�h<�B��@�A]����
/^~��'��ٮa} �h\�����&�P��D i
$��(�D�4G�hS�ή0J�&��J`��~H:�pw��J�rf��8�*�>�'��,*��@舏���s�xd<�0Ω)����+Uq�WMӽ�ܪ89��H#�9�?Y���>-,X�e�M�L���*YP�����Ynh�0�c�u@�h�d�+UϚ����0���� ��m�A�Y�U��"g���o�%~�BA�K��������D��tus3W��X\��O�Ki�Y,PU��%j׷�����ӎ�K*���I��(ی�T�Ͷ�lo��4K���~�=�K�?��*���c� �DB%E�T����n�VQ%�K�^@:E�DriP��EZ�����y�#,�����w�̴��0���$.��|֮l;ځ���e�����Ǽ�ԏ�+҂��u=��g���:/�;�(�t�Q_0���R���z���ME��mCCq���i��<�����E���I���E����ʊ�ү���׸�Y�o|Yܰ�C)��]��6OO{�p�<���tՁr	��<���F����Ys�����<@�B~e��c�*��0P����h��~�<��_�1"v��uD���il���2�����q�F������j�8T�-ܾVXV��h��Rs>�Gk���̔Q��t��0/G�iO�vs������,l�И�ѡ�Osm�Q6�c� O�
�눛�؟�#�a�m+9���׹�=��Y[Z�P��ȅTtZ���{��]�I'((�m������S�����,��$�m�CBg��uH1��o���`�ײj�{�۩`�r�Z�e�6���ܔo���f�|��2ѷ;jjj�s)��N����=*O\Ěz�����\�`:z" (�]g�P���׀Ic�/����g�]���=��-���
eܹ����:���V��K1���oG�"Z	�0GGjD���2M�B��oD\f��H}�b���P�̻�Ys�����q'���\/��Xn���n�W�_WB�������	'�bEa����}�rR���a������0m��3Rs���o��X��p?�G3�p�Up �++�ş�M�[���[1-�a?��,����������������P>q���2���P�&��95sE�x`K�j?�����ُ������emm1��>M���MD�����b|
�-��]��w#�Ε�t|�,</���<����U);�|V�y�f�� ����e��.[�h)HT�RGlc�9ؕcaL!��"<�UT8��=#-��NqwBL�l�o#�0:ha��t�f�x����l(�DȖ�*�3�����Wfg_I>�?v������U6)IzSܶJ���	^�:s��������h�L'�ώ}�����j��b�<��zl�n��R<�3��Ɣ��t��S��jQ���sL�@��3��՟���W|BMI)x~�֠)��-�?v����ʬ0�)A�0�&r������I���1.i���������sN��t]�8����K�!c�[��#���6��e�r��&������3ĝO6vvJp��~��[��b�3o�v�
���j�툅�AYy��l����8�Khy���t����{�V��ƞ������;����x[SSHIIɻ���(*�͒���=�)�9W���	�sFje�cq�c�L�&P]��3?��6/t�8=
O��ģ&�I�<��ׇ�����_��o{+�PKv�a�R$��%@Q-I�{���6������]�T��u�����,I�s�5�c���e�Ԥ�B#�N�[&e+r����~�8cL��cbo���mo�;���������Q�zŮ�ŝ��HM�2v�
I04r�W#:Ú�L<=u����a�����qN:�喕E��;����Z���C{j/c,��o�TW���r�}����7��K���W<��I�6u62��646N.��F\�ț�!�ݣ�Ө�L��(��ɋ!
/|T�<��U<�ozq��a<�cXR[ו�can��2�=ˈw��|���4*��5~	hd�9��L5�i�ݯ�A�"�B5�.�����^��.Pbn4-m�^u�|�,y��!+��v���C�eZ���&Oڽ���=������x�G����{%v���v���\6�"��~����_��n����)�<F�*�c�f�Ӕ�yo�g_Cn!���wY�gM��������z�Ь���c9��`fz��X�8���2)<�X����Ai�K_H,���T��	�(�5��m�����>�-�E[LA��ED�a.�� �muH�����l��&x�̺��	
C��������j�\U��c���bt�C��R���n>B� ��W�\Q)�@7�)���^�ݜ7�]�	�6v	�f�X���T���*Z^v@N�x�<�cÆ#���t��e��X��r���U6���3֜R����'����S4��M��]Q�\	w�vI�V�wЍ��q��I[q�%�~B�jr���7�]K��1������=����f�jg�B"#Qw|r����͐�/��s��,���m���g������힒���9��F���h�Ξ�Ԫu	
�w�T�N@ԁ��[d/�/luF��ߛ4�c?3`�l�������Gd&qo�c��n��Z*+l߀aQ���i#��^�����We��,[�����z@���7&���fA�ɱ{+���
ov����J�W���\�&���pOQ��?���n��Y�i�R���D��a)�5�(�� ���ی�R��ʴ���=VV�ޣc*�A3r.���G=ϓ����t���9A�?5V�[r�i  Ԛ��AbĀ�+�dd�eƛ�8l,�bDʪ:8(#�ݭ�ey�Ihm��>#�Բ2M|�G��RY	F')�^4+��Q��.��2�J�&�z�Wh7�����c'����z�ڿ�b4��-�G��6o,���(sjk�QB۶�1�I�� #e�V��t�xe�o+rv����./-�R����sv{J���`��;Qc�R.��*��,4���(툞��<ԙ-F��\�X��"5����8����@��|�k�`�#���F�yu���δ8f�=;33$-��#lz�7d��l��vw&��MuIRLaC}{����ΎuD���0���g?M���|�i�������������QN�Zݨ\��ܯ�,��5"�(�֋�&�Y<^�У���	)������xٹ�4������'/l�c������Sl'�i��yrr�y�q�����¢"T�6555vw��>w3����?�;��U�������w��1��ev�@��<�zZ�i@``r�5A�/���m�c�u��}QTZj�o�l�
�H�P�P�h�����Xf�g��R�����}7f�3�eb4��{���L��o�C�,e�A�x�0G5}�]g�C�?ߞ��E,�q�x�۔[D$��D��F��\���=u���v�"��;ZN������4���K>5�G{�b������o�����2\镾=�����e��(t�Ǽ�w7Z�\����͛f�A��5��n������̏�X3�<~c}WC#RUU�Q����-�lx;�U��\j=�\���8����r2�v'�����8�Oz���Z^�O��۪Z�+߰���~�䛺���������*��+��	F��E�5��>͜u�[f�)&����@��RQ����QS^i��d�5O��|TYQ�񝁴���c�_��;���	��ѳ��U�dj�VXX���������L�ի<zs��"#�
8?𽩣O�<�ߚ������-��̗����"�	&5�� ;�73K�2ibb����,�R�f`�({����[��Cp�U���"�!��TSm�齽�t�.��d�ȤYx�F}����Bu��I�C�n��*)a�ïNb���[�s ]f`N&�4����2q���p\ ?c�T�r�f�eq$��[���")�Zͼw�5sAqE������wb��L��l�3��k�Ȯ�n�;/��0l8�8�me�|��R�\(����$$$>[?�� �BF�'Z�to�����x��QK�ַ$l*�������$>~6��ӓ���S$/����A����dWx�V ���W�M;}����?��j�UL:� O��x_��V��&U��$TuJmzwG��~�����Q$	j�t����c���~B�Ǵ������e���]�
�G�.=��}y�r
:�揉pp����KI*�T�o�ʜ��}tXZ�K
ڦ���Z�Ś�<z�?�؏ .���=
�����CJXl=��5��� 
A�m[��A�2�622�ŉ�皂�\D��B��-,,xʮk���O�u�U�]mX����9V��)#�VH�1�ɡU�e�g{��a7$�g�͈��Eaa�0V���0�y��gϢ�ͳU�ɇ��s���9M|�'^ԃ�	���sC��q��{�W��>O�D���$K1xu/m�������(x��w��f�.�������5W�ޭ�q�bHF�и�J����r��ױ���؝]\b�ڗ��8�����[�>wt�N�!A淉�q����UnC7
�-�Vg�@R��]n��	�7����,��]b<��HUY9)Y*�"FX�/O�k'��A������d�zcD�Q����u���ǜ`�RIW��ݯISJ��x-X���s�˩�����U��	����Լ�ٱN#��o���Z��mm�W�ၔU�X3��h\b;�_ �U��Q�M$�9ݓP�?)i'�^�}���f/����ZL�]�b`о}pl��C�`����Ȍ�!q{�z0�}��i-��j�f�)�Ú�����W�c�2AS�y$2�'g�/2��X�v5g4+;}I*��Z���zÞ���	pp�q�Lp�69 �د�%s�7��}m��R�د��Ƶ@[����m�Ģ�|�śqk#Un[ŷ�w�#k�Kk�8�44,[�8�W\�ml� 1VA6Ϡ��\�@�x���uT<��F�d�T�}����q>|>.Zd;*��p9�_
SiX�|4��+�s�SANw��$�ߟ]X(v�J�+Ӊ�Va& �WUS+�g+mw{�'Y��0�s�I��v��hK0������=�ꑈ�Z�'1��Ͳa�] >�p�@��Դ��o<5ϞnK]�e�Ы��C��������r5Z�d����U/�#��;�_]��kkޑtW��H���Zts"lko��s��#�\�O՟+��;G?�,L6��%*�Dp8�4�-���ZXY91�<>�m��f�l�e[,�қ�����.?���x2\�j�K	**���.n��Z4D�/I>���t����im�<U}}���!閣E��k�0��7j��e	��=��-y��*7�y"l_����Tk�$QF�%E������&�����@�mO1�j��~q$eF~�i:�+�㑸܍�_6�J�D0������<FO��'�CL�z�hA��&�.������:z��"g�����L��c�Tk�Q)cj��1�2
r2<�[�3�����W�K��z4�Hݤ��4p)3�@�Տ���i{�ؒX\O���sa�u�7TOO��j˛���1P�,7;�;U�������1����`$&b?��S����ۮM�)^��yRE\�˪���ޭ[Og�	��ώ-]�Q��4V�kg���-(�kje�ǲ�jc�~���A�X�@�Hq��u��c��xC��#�ZK�єR@pW����,i�6N|�~q��Ѧ�@��o�Я_�����DyVC3��ں��`.��6����u�����3����?랇ř�~P���4���X7�4����no�'k�����@˯��	s���S���Y�߾��;L*�Gfe{_��r^�c�;�=(�G��R�����;�o�&�T�]��>M<�O�$tn(�(eZ�3�*6Ĩ�1r��m�tt�?�1ou�	ƋyH�8;�iRs~>�-g�)�Q~�/>� *&$���>k�dfN+�>!��Ͳ,�}��>jٸAhٙ"�74��XD��%�7O��JBE����?к��⛫�����K�+��r劣��Hc�^>*�X[[��cRCM�B҈ʳ���/h�dxʤ.�<�Y!���o���kh�"�]$�����朡�TȺ!A��+��k��Wk�c�K�K�+T`c3�掝8�eg1}��4 d��Y���(]��g=`l<�9߰��Q�E�cH��!���gu��Ĭ��W��ӱ��� ���R����ɒ����><h�x��\'Z�0T�N�Pi�K���܍!��Y55#�G�?���s�JxB�|,���eH��38�G'���v�߿�TB���G��k~U<:�|��kۥe���JГ��7���)��Go;ma��֭}re��}�븘��լ�ޛ��a����&d��y����ï���B&�nS)�����:���EO��������q�ؓ�:ુC�Qge���*EŪX�5�T���0���0A�O,�m�zp�p�YK1T,�=
9ޫ�EҠ��C�v���+��%a�1�<nl݇DjHK�2���lH�fw���[\Ă�0��kؗ�#�����,m&7�7b�I�V�Z��K�7��]�qV�JQ�>5��{��A����V�HkZ�~�s����Ou[�06|�MXH���{��_��OMx�y�!�	q�dA���7٥��n^�w1QW�P/k�'**ʧz��.����"))��;T�Q"����v��Am�t�őj���Y���*�p
^�޲�{��o�L7�I�#�2EA���[`�����J���KWv����(y������\h�`�T/�b��N�~q%���S\z��O�����@��O|���m6b�$W&u��"����]L�A"�=btG9�E�d �.��"������M�?�U p�#_���^�ܜ��fH�k�C'HHt=f�d@�Y;I,����@�^�:��5�`t{�֠]|��`�XM_?/R�]����۳337"����V��;o�@�ϓ�[���f0G��;�V2��w�n:N����f9H�]��{b2�6������&�$�<~0;$$�N�A�������#qj�
v�v�+�����r��au�������7�YV��Y����]b=�������z?��^m�n�
;ם}�8r�H��'�?�b]̌�V�5���ɏ��W����4Ќ�1�b@�6:��	κ]|�c��cߣ�2��,,��H*�izT]]�V.w���E����[�,�����n>\�&W���H�Dc��Cρ�E��oċ����q�� ����bȫ�"��%��>��&�7��ïh8A������<�$�����a��MO���M�����<�����ih#�bUJ�6؛4����:��Br7;ہ�,��a�r���	�~Y;55�O���%���ѿ��H��(��}{{!M�@��,�A���T�����uP����3W�*����������&�d��h~|R�5�ݠo��/��C�l�f��0|�=NШ��ᝋ��mlwZy_sZ���*9P1� -ւ��n
cu^�u���d�G��r��ɒ��E�]<Fe��@.l�	�'w48��D��S����Tma�&&��MRQ�Rg�XZπ�!�%��ǄYʶw������
~�ȡ�(ݶC��5d�|$��.D 6A�C>���@�M_��6h#P�&L�UUC�T�C�w��E�x���'!���u��q���ֆ� ���{hh^���)e9�7����}}
�|2�,�	R@@}[ܨT� �y�h$>��5����	H9��
�����-LHDDZh(%mv��#D�e�g��:"oW{ �վQ����O���近G >�n�S;L��ch���*��wP�2�@�G(DT�
䀋�t11I-�*3v"��>�`�ӧ'!����f�� j��s5���2�O�Y��u=S������h5z��>�����P�;MA]����
?EM��{�3B)3Z̫�J�ȈϾL���_Q��?�&8��.
vJL�e�K�G��^��=�I=�k�n�KUK�	�q�5�WX:oZhx�1�U�,x�sy�E!��׶.%�e�����0�6-�$/���6��P�A	�����v�4t�A_�a�*��ش2��Q���ª��$��A���õ*��C�|j�ddd����ՍH�/�?�;�ޭ�aa�F�����U����0�/�lԵ#�~���v/�8W�Sz���� y{LV��(����	H?JYII��ʠ���mۚ��
g\�qY���n�]kq�G�!F�>�f;w3�qP�F�c�b|(P�-�RE����B(�]5zA}��'�ugy�L��a�j��#7=c�m�WV"E�-8=��V?�����&�7T
�Q��ܒW=���a6����ȩ�+%�鑜���Ⲳ�bx���No��s�l��B1V��h�?���׳k�׽���^�07b=�\���kH12��&�u��c�W2]��-�w�dK�ï$R�`�#��a|D�,y�l��z���"//���s�S�.���Iru ��?�M%P����f~��-�����)2j$������^,lOg���r�"��a���03q���F�XP�ϩ���g�48=���޶�jl��U�g���H�@!�ǯG���:g���&�O{M^1�7^�����,dV|�U���BV�3N�m1��:���u}U{��d�+y�U}���^]3�:�pf�KBW���M�2�s����]]F(�*O�:�QT�l�u �Q	u��M��0(6�`�^�mOM�"��C_D���A*��U��y��щ{���7��]Lk�I�9S$uPpw�W)>��N�;�<c�݋��]J �H�'�9������ˠ�+#g۹�)P홊�2��z�y�%�A#M�BMk���xC�����\O�b���c�l������p�����L�kG^y��㋰Ʈ�4n�z��EL>�t,) �$�]���m�����^$�R��H�wyⱢ��V+y㧲6gI	���6��ߗ��~�ZR��s�q��2��<B���o��D�5ۭjD9������R�ȟ1���e�Cm@D&��]���Ў-��1<��{��}�,2|���3������D�)XG��]b��ø�����F�62߿�T��F��O�����􅪅�/u���l*1�E�(:��K$8����N47����)�v�{���n��'��뮫՘�El�I�y�%��(���Y��Rq6��<޵H�G�,����-�������1��!i��O���}Çl@�j�C���|�}���rG��)�,�2���ÆdbfS��9�];�&'S��P���R���ģ��TT}��&�U����׮�,����uE=G:�-9� ���
R�k:%�3�ttt%9�K�uw�;��kG���W[T���(����*�+���MϮ1�ʜ��-����҇{�¯2��\������ȃżC����| �O�&��D�	�$}=�sC(d7n���e?DЇN�^�j��#$��hx�
�kgs������̇��-�̎C���l�!���3.i������>F�%���Z�׿��3����ѕ]�xz3��C% ��DSXޤ����^	�R¼lo��x��D���ɳKJ�Q�XG�1�VR���4X�Z\cjzz�CRO�G������v���-�֎� �|��qJ�QWa6�=�������4���X���Ħ�_�V��q+�E��k��,Iz�))a�ԲfģKWد]�Ӗ���ةspo�&lo���r���������&rYN�ѦD�������ؓb ]4⦦vW��f�Nw���|_ܐ���!�&/�A���!��K��g\ބ����k���$!�)�J|�T@ts`|)$v)S(�A�.d��EN5��Nj"�נ�D��P���[?�A��P�8n_D���ϣy�X�<�j�F~S�����=O���wuuѵkiq�Z�|�aucuH��9V���h�{�1Tink���ݦkg�r�r���&Ĕ��C����͇F�I	�;�虳�˩fo,l�ֽV�^��� �2�ځ�9ɪ���s�#�ϲ;�~Pn�B�ɉ����`��u(���w��"���0j ��}��X�W��Dy�����|�PXG�ȱ���y�f��r��t�x�|ޅ%.�y�ł�̘������bcem\Z��H���(t[1m�<��cO�:�sU,*,-�},�ש&�@F����ܷ4��&�X*���<t�آHgum�ajm�ڍC�����#��=��X�ϱ|��^]�R��iuK��s���cP�ib-�����z�pIN�U?W2٫J�e#�䂝�k��h����ڰG�ڦWf���wg������g����-�`��ܜ��wbna3j��{vi����ƶQB+ݛ���ވ�� r9l���������֦������'''�U+�
�bx[������d���/����H�����u�2����\����C�6�
���0;���a��e*��_����<�#"F���z�w�ė��S��c��SuDN)u��fo�p@>*..������Nlڞ�{�|����Ҏ���EJ���H}�!
��R����ɣ#�ns{��h��w���Ŷ2$��+�t����V��&��JF��9?�̮�<���87"��mP�yֽ-mmΫӯ�*��=*�g�'K
��
�Q����:*?A���c�_X��QR�|�3�Cg��ϟ�AS������3A�%ov\�qs��$������A����d�l�f"�J��s|����D�OsG�BD�.> �m(lf�������ܽ���cḿ)���N+쒃��[<u%P
%��̭�R�w�K��Z�Jm��$0���M%�=}i�1t��Z���δ86LI�F�m!�	(\[�Y��lJ�t���V�yΠ����sssׯ_o�X3k����R�ib<-�E-"�'���Ǌ�x����]�i�v����	���mݮt%���;X�*�b8��|U
�����Q/��LL�Ɨ���o���â+(ZW�H���(�|f�{r͠&�K��M���^���:퀇���%kO��T�ѱ�*>B'�$������bG:��eoNAfL]ff&gC{Eee�㴢��]\ ��_9���
��p��d�(,NMQ1�xX�#.�(��%� Uw����P�*�u����6��0��sӡ�Y ��<�q�*rz��o@��,��W�M}+�ڰh��i�Nގ��W�i���+��^�-����:�����,��G�Cyy�U������?��b<D�9jtm���<����&GЂ�m�A���_W=�
ʛ��De�m�ୁ���RI����$�����4-��݃��9K��ؼ����Z�S��כ��8Q���)s��R������2Qv�)Į���Y'��k�כ����.I���/ϚѫtQ�X��H<>�mmD��[j��������������E'M����Ɠ�.g�O�\.
z��Y�x��4K��M��o���:X펌跰2�V���Y�ۚ��@?�-s �zK��g��m��umD_{c��9\D���O���f���UT��0����3��׿�p���������6i�W�fR~2�p�KM�B�^��C�� ��7�kJ���޺�OCC�~�z�u5Ȍ���V#U���/f���tp��w⬿�>1��}�@�_�OC�ʅ�jzz�Wi?�Q�y���}~��i'��$x.7=��m�"��LNNnrc��������� v7ޕ�=��a�»������3P���u��ug���q��ܾ.�5^y�%��V}vK�������xY�ŗ@��Õإ@`�p������bܨh_�]�0!:��|��I޸�7��f��A����A�a�MwB��/ع����v=�)��7���Ϗ��.Z���N������Ac��7�e៿s��{w��o�-6=)��&A�ƈG�:/̔M���l�\eK7t�\��BK=:�9�ds�{�_�ԙ3s��������6�cbb�b~NMk��&�pŋ�N��{�J���Ǭ-�C)��<�+580�;J�g&9xU�?5V�о��͡�/���Y`@g:��L/���f��}_�+?�Wڥ2�J˪R�����7���9�[g��\��a*��ՏL�����2��yN��G[���̌�B�Eii~��� �y-ޙ~��YqFu������Ig�6�Ѿ� %�**6��R?����`�e���Օ�����8ѵn�s�6q�Ѿ�+����>����4��}Fz�|�J�^���ڭ�Ze�N�p�lW:����c�:��\��F�=t�}8�]�u�Y���.��׌�>7��[:R�:�/��.�������g�K{"�[{;vZ|�m�mt���E�����(����~��`���qVNě[bm߾�O�Uwc��	��{��b��!���,efff:�ΥA����v�曙���*Gwb�Bvx-{g�
�|kFƗ�zw���F:�u�������� �����NFG�%Q���NG� �n�{%v4��v���o�/���e�4���Օh�D�7��3Ef�3����H����݆{��rdm���4��4`s�A]=BVNn��������:�稩`$�ց.���TY�ݑ\[[�_��҆I�TIG��}���
��f��+]�q� ���N���LZ"��M,,-�F�=�}!�rn.V�,I�
���F����X�d�/�M,�b�{s���jG1��wcgc� G�J��g*��]O4��'�����XXh��EK,�}9ō���`�V{��xԠ��������bu"L�\�~��?:$���^|Nv�ΗHPLX��ߦ[�f����W=�����5��Y���5�)J�Y�M��l(��b��ǧ��Xl�B,�`����/���z-�g+�T�����|��[,Q	쬊�I�T{���F�"�R�->>�T����/���>�4���NIKcѫvW{z󦞞	�����̣)Mү_��U���7@1�ħ8��k��Ҧ������ u����VW3jk����{��$�?t$KY�G(%�ݠ�oő�ɋ"�zBd���NW>{vXt��Bl�aj|'���ay�e��YS��ٷ�� �%B��Z󝛛;<""0jݘ��퀺u���ׯU55����������9obV�^�a��f=
r�C/�x�ߴ�����n����sb<���w�c�SQ	.U�N�7�g�]G{��6���Lh���ӧ�l}�3p 1��.��c���;�!���#����뾻���N��<�YS��X������
��Pr:���N�K�jjj`&�y���;�n97����G�=e0���lll�� `��g~\����oacS��'0)5����(N#�p5W.����A�i<|�w�-AT-�2�	���E�/�=�fu�	x�9O� ����P�}t�R�F%��ƶ���l�6�[�eLl�3�K�	㭅�jKl���J�D-{�(9���������G��Ws������WI�gii�Xp.���P��GO�߹���'��Z]]�GL��^^^�:�
vJJ��6��d|��S:"E�y�h����SDѨ�:�.kn$O�:>x"bO�Ī#9X̂��V-I�b��h] 3�X�i��Y�%r�I�Kv��y3��ƦW|E\8u�b%8��.P����q�[[[��YA������_=��	!!�ͮ-롓\1���?�|A���ķ�<�}ţD��o��/����e��p�=00l�����Q�R�b����k���gFm3��#?/\%�&�,���N���]Ď��ُ7F�Sm�h{�.C!�Џ1�\;�����[���]%�#�HtvuNb{{�����e�d��[fc��t�����{IN�z�B-[�Ƨ�����
��}"D*�����3YEE�	�4�����=�t�C��� x�ut�TU'�K����e�'����WB7��9����:	�ekD�]&)ﶶ܏~����g	�!�i�C�F8T�h�í����yz%�h� �KԱamyQ������Tx(��[�n��qJ�����H���Q�!]!��'�d����ߊ���Q{Th���TZEgggx=GGԃmq����hy��tJ:6
f�aR�����#��9���btU��=9���k��X�'�K��Y�y�ή��g�Kٕ�:���|z����R+Ǯ4�L4�;�C�������?���>>���0U�$����CC9��.�%dXD�׿����N�P�vY+z��������'K@P%���
1w��2�`�8P֨�`i��������f0PVN�'��1���7�԰V�HhҞ(���U�ZM]}���R��XmvU�������g3lbj�b��W�§�փ|(�{Z�h�f��?晲Ā��=T>�u�dyסj���/d�]�_��B�paa!�꥘+>	���k�y�i�/�C� �f)����h�Az��2zKB�WgE[���T��;��(s���nO����]X�|��;�c���|�k�]��}�F�Z�&�ɩ�
͎����<Ro���m(�[3O$9��m�;#%�|�T'�]B=(vm���7Lk�Ck����/ c��n�]�|y�ZAʉ�@�/5��l�+� x�.Y��oU�n��|�v���Cem��� 7���42<d���Б���� o�EHp2���K�����@7��u��3�}{4��U5�Q�����)DW��
�'��]����ֹ���Y#�'�ۊG\+J��}J�d 
<��y��#<7n<`ڟh
������U��E�$��/���Z�?x0MO�K��	��^%&���j��d��ի���Jq+��o��{)&��nmo��C�	�@�G3��e�.��먲���h.B.�5>!�oD�t�0��q���7|w�HYeȫyG�{�ރ�^G��@�gٷ�����m����,_�j���&��
(�씔/7��������;M��ӴT�X1���^j���I�q��AQ�\�ڑGdK�d���v&�Y�29eH�߬˄�"�z�W'���h��8O/??n'q��"e�u�M�]��."WNx������|Ƅ4N3鹮���{����"��K(F�G]	�T��bh�sܢ��&����1�b$�(y�4������*t��|;�剥;�?ٰ(ݗ�d��a
?I��1�Z��Z����i��_P7GZ˫������f�d��b�e?_�7Lf}�ω��e�cygs�He�����0�[=��%t*���[ͶW�U`�)�A�bNl��f�	j**a�\�/��?5Fy�� `��� �Qd�{Nx"�j����*�(�w4�����eZZڞ�·�+�V�l���}/�H;�#�0q��Y�^*Y2�b�������$��)2��ͅ�����S�Ut�#�sHL�9���t�$�59�B�?3iл�.�ؙ~|mc糋�OcU������{���и���+H�t��|v�>s�����{��moKk��v�d��	������nS�.�HKt)��"��_�U)��ϥ��-TvR��,%/�ە���]�}�HUM��M��㥼���g���]Xs_܊�����6���T�Тd�(}�5&�뛳W�����E�8�Zm�ʑ}��Mo�te�2�+dnnn�[Ei�|:�Ne�c�����l�U�Ŏ��%�I��n-M���G��G���ɡ[��!��������?H�1��݊(�h
���LB�dm5)y'�93eI3%Azy���oJ��Klj��-��y'��``gVp�<�u�����h8�:򣣣��~Ł\�[�v��ǡ_է���Ȭ��h���ҟ:>KOK�-�}�@�����Pf9RU��5֭Z��D���fY�r\���%%���ݧ�]���t`Q�{�D+̓�`im�>�~���`)�.��v8����5�qf]���<<3��a���@��*8>��
g�*��
?Kn� ��������s��� ������l���n���fG�5�n��:/�vM^��Nmk [�f�;�aamͫ�|[ ���/�0�R700���Ǐ�^?��)��t��Id[�i�T&�r|�]^^�	����ӓ:Ĺf�_PxiY�7��C��0��>��=N����ս�U��HgMx���G�А.�v�4lgk4�^{�,0����4�G �4ܦ�M���N%�-�K�7�pss���h3�"�G|r��$%\k����-�4
MC7�|�^\T��6��<�b�(�w��G��<��#��e^�䊶��U��
a�'΢�II��=sj`�*�t ���q_���ɽ�uK�`�jwlצbm�~���c��M��+�k��)�Dsm����
��� ��A����	���)�H��E��`ɗp�Z�+��q����XetkS�|l��X jL*��ÖUTl����RvǣX���h��^�%����dB,�}��@Q[��-�[b�	,{b#o.�S�'�	��L�i-�
ff�HF�c���cY������I{36&f�W��|{}�uX7������FE��f�:"U��WH�Z]�G�g�#M!5vMz�3Q��E���5Eǌ��Ȅ�G�^�QG[� "O�j<�7��ͮ��G[�;�چ5�H���:M�� Ш��b{�5�`n��� ��*D:(I�ƶ��mt0�;eF���3���z���;�;~fffT�+�A��I�J���A[ZK�D^ˈ�oޠFA�N�t�X�����v��E�Ӽe�Q�h%0�c�qp-Z���C���*��D�(����z��c���;�t5��нV��~��l÷��n����P��yxD�Eo��}a����p*�@yx����&A]��e޻hБ��r�:á�r�ę���>'s��%��c�8��q�N��@�֣5z��$w񣎋��J,���͵{p0{w{�t�@���瑖*��PڀnW�\��'��c��4�:�%�4�ЉJA����� ��&w�F2R=��x���o���ϙ?0�y-��,�""� l9���xyyiZ|�JM�_�3��ǣ~������v���8��uj���U�a�D*�ET�M���|��&0H�mZ�����&��n��+���d矙�P"$/n����SQR
vww?u�hwWWrPP�����~���h1�@���䦧�wōQ�Z|��AG�ׯ_h녅��!��Ϣ�k�J����d���żݫ
��:���7t�-}=�/�(2G}����tѭZky��W�b�X.��:�%��y�����yP���zi-X���iޕf��?��k�����/�-�u��m�=)HI��߄mmm�X�}˄�f�Jݪ�A`�ٕo�z�GJ�l�����J���P�mKCG0��]뚼����R�!�,(sm�<B!rr���&oO����"#1���9�f˓/c4��N�L�zmgN�=�C��Syn�0�S[m:sM7#=�{���>~t����p{kk�L�C�@t�$vif����5�P�{`�B����0v��������U��D�S�%1�R�fff-���u�Dc�U�v///4ѳ���]��6ף��6�|����r��4jv�$���>�^��D�hvnnAAAY%�ڵQ��ō�����/S��na1�'�ihD�b&��^��]3 m�!���IHHx~9���W�UG��%��015m�7\�-Y��>x�`�7��(2RR�y�a�Gh1ry��9w�˟]oT�Ș�]ܸ��:�+��4�qH|�W�?�B/[*<sb��)�ᒧ<����۽Ҷ�pH�^mb;J�2P��N`����WZZZ�qUOx�! [u�S��$Yݦ8}ɦ�Q�������� -Y��}yo�x�ӿ��7�ʊH����bq�����#f�N
���
j
����U������>J)���☃��c�P,����*D��^y���F^�5�I��ˮ�'�P���c���)���3E�����v�����K���cގ�D�fx������2���4��9���v��!�5
�8����1z�|�X�Ec��& ��%�����-�X����S]BTC��I�:����%��Ss�����5�v����t%WP�^��a��҉��1z_��jɴ}��������@*775�s`jjF�����'�sCF�n��\�e���!�x���A��]~�!��,�R���="
z'���η;̤��u �			����NCOb���]?U�%��44H��	��Ul>ԉJ���������(�-.,gR��GO&������G`��>�������G���:;�����C���]]zM��\�9�B� i�S� ? j���Q;��_��knn�m���P�щ�w����7��r}���TrJ)%[�҂l���c+�$d��cg0T��+�e;Q��a�CB�e,��e�ih���~�������ߟ_��9�����گ�u���<x���j X�d��G^���v����A����X����}M@gcv~��(�����碬#k����je&&&��>�e y��dY���,��4}#�>�
[�������I��&1c4�p�[�'
U���`|W�i���^Q'�2~4����_eL�=V��z0�\�7�*�XRW��є�N5�H5M���V̊Tބ
?tŢd��;��|���8���a'�3K��{�G4%7��B̺@D二��T��"��+�y�"h  �ShQt�7�ʉ�X[q�_**d�w��A1�0�_@�g췻F���� �Cߪɳ����8���ѝ�@�?�n��~�z�ȭN(P{�}���<�;��/����$��ʰ����1�I��V���f��m��Ƴ�|�N����������9�A|�Y��K��O���Q��.��m��Ł4B~"���������������N�=h��7�;�/��3�����O�HA��� ��#�]�شri��P�5�i�*�� �#j�Mڪ�3�=WN�}S�J�2u
��q�$	���̌K��͗��+��V���+���\�` ���r�;�Q�������"B
dD�4v�KA}�P	@�ni������������i�j8�P>־gb�ϙ��Wb��� �����~���������N�e[~"�(��Z��тY3�q�ؾ&|%�����~/hOk���1�ù���8}�ׯ@�<%ǅ���x����*t��~�F �d��7?��u{�����0X���v�f�H�n��'��>�:`F�� �`:����,���4}.e5�ٞ�{~Z>�����C{��������`���8W���� 91ӪL���b�x~�^FY����%$:���,����|#�J^�D��fR&۟�<���u��Ι?0:�ݖ_������tF|sT�kh��\��A^��=󈲽��?��fdB]�t;���M�<�P#դ��&���i֠���>R���q���1����i
d�MR�"�T3��HLO�<��v�w�0�Ӏ���>�=xT�s�088H�~	��D&�}4rO�����2Ȟ�>����o�F&I������pAHl�^R��o�u�Z�\�'�ގ�) ?C�Zn� MPo�@�m�����cS�s�\P��y���-���P2��j��ݲ�N�O����k鰝��v��emCR�"��P`��b/}��0>������@qv1w[��9F�O���~o�����%	?
�O���A��uws����Z��|��@�4	�3/!�I�·��T�N����;Q�&��nF:��sKK���]r������ �x�s[[LӘ60�#?r'� ��LMA�B����{ol�m���4�a�{�=9������$t�����~�h����_FrX?�C���S������>��G����u�%¼~Ѣ;��vw���y%���8>�=�N-9�SZT°���C�7�R��Ȯ�|��h��j\}��z���>����͘�׸�
;/<���H�I�-�(|&3�f�-��V��-�Vv߳ո��	V�̘z'��=���y�`�·�����#���H�駩R+��`,�Q�{�A��%�3Ie�X�y����MS���+F�x<�}�����ƁkWM�4��\n"�k��Z�h��QׯQ�`bS��+	F*�+p�x��Z�?���?Z�A���H��M�Q�J�X�*�b/
��nb�[W����zE�0�V=�F���������ARCV,v�oD1��Y�H�#a��G1]��
YK^Ji�j#������_�1?�U��%�U��O)��z=�I�I[.`�}a�#`^�ךaJǽ��Mn��ϩ��uO
�*0�[�����z`s����E5�:����Р:~���uO��_})��L���ǒ�݆h(�^-��f�	��Z������gw�Ag�����k?�޲ί�X��7÷~ċ�_&�,V���"ی���{?YH,尒z���S1|s&A3��������ei*���) �.s��h;N�"x���ӭ^�N�P[���7��o���KZT YL����:���(�V�BT���WE��z�(�Γ_���y�o�~�XT�E�UY//�AG)�W�a�io�h���dU���B��7+�t�Gu�ե��H�e�3�͵u \+��?��`�֏}����u��=�au5�l	^!���3��a\ډ�������ha��oo5n4�@�
g�� �N6GV�r���K�}"�3sV�f�A\�g�a�Q��H�=dܽ���P0Q츁"�f��V�=n�a�Lz�@�n�'�C�(L��=+��"Dv�x���vSS�+�Td�ujbÝj���/�'���+dg�����?[��AG���˥w�JgC5������IJ��\�j� �+	.I�w�>qS?ǜx�ӒSQ���-	��.n
݄'#�X��({W�N��몳�E4��î<��:)�3P�H��%�-6�[x���[�"����������H�
��2�����2F�5����KO�)^���1�\�a�縢�9�O$/�����O�s�ݸ�M(9��F��:��z�=�x�C~-e��S�6��y�_�舡=e�D��%�964����٦��9I�0���.�����J>�4-��a:��Dd��dB���<ϴ�+V�,<A�I��I�$��\5���M�=� >3P��;@�,�ǎ�t�8(��[��bS,�r�s�|���o�k��6Bk�	��_����_�~���7���5��P�j��/��k"Z���ò����
��g����;�ad��MY3r?bF��m����lb�St�	���AA�J��2jK�qϒ�ױi�I��G����	���vu����4�ڝӗ�c��4Χ:�[+�T�Y������7"}�O6/�s:�ɥ�Z0x�Q5��ۯ�'<K:�"}�'%o�8��d�#�G}"�7ʚ�`���{Wk�~�:*��8е[�_��2Ο����(�$)kڬ*]��2�Mc�r"4XP뭭�윪?��W��&�ýd�^������^[��$M�C�$����y��QOa4Y�L�{9���~�>����u'�";[�)���r@�{?0��]�>X^&�m���W�y���O����-��m�~��*JG��M��'��1���%^��α���u�:_�(�^uA҅Ԁ�u��ن�E^��7Tv���(��pCJ8�9���r�%g�����D���1[D6�Ce��+���OOg�"ʆ�p7�r�?u`��2��a�	�ϊ;:���g������f9~Ӧnc�_�cY%	s��V�r�rڥ!�Ǌ�jjj���Ńg����@o뭞�g"\� ��"-k;����춈T���a����N�ju<W��݃t�xp����ͳW� iCD�Y=dTc�q��Ey���tm��nkqH�O�ؿ���:{ pUF'=���T���Tn��9%��[�LZm��,�	�!���՘��/����
Q�R���8�&AR��X�ܱ��Jq�����Հ	H1G���M�\XU�O҃�I5��F+�`o@Lx�@��?hh��Y\n�nNA���V�k�	�-kz�����O��w?!���?Q4=q=�$S-��v��`Aw�٨�� �6{ޡ{p�TS��m`an`�~4���R��]���*�2���Wd���T����զ�:������m�3}?���_/� ص�{G���=1�������VR���l�4�D�M��y+�VS>���5M�|��jV�����b�O��=< �e�kC�qE���V�B4e}=�����z�7��υ65N�i�WB̈́s-Eӿ�t��"+NxP�DP��o�o�;�i��ۊ�Z�n��*`�Lwb $�%�:�/� ��d�Ng��j'��,��m#�e�A9�͸g�5�{�VU�����J�yEx�7:��1� ��r���9')L���*&��@� ���po��н�E�{�Z5�Fv%fV�����Г�������M�����c[�OQ��v�`<H�����8E�k䣫�c�y�6�(> ,�
L�NAE��[���Q�y_����O��6���PWg�\�yc���9�H��O4=��V��R����W-��R
��4(���G@�/|� �7B8�@A���%Z
.�)�3��&�)�4�Z$�����z��e��isj� ]�<�{�p�P�>�aMco�����#*�riV��ke���q	��&� t���^�VHI�N9J�81�"<�K��K/-�lo�V �R|��9�<���M?uEYm[����DH��>������}���:CQ��+׬��3�& >
��)�{�:��S�@�r{�F��aZ���2��+4����}���	g�t�1��ʧ2���^Zs�tgOsP�>o�N(F˘�v��ZO���H�'p����YT�V����C���.hm���s�N�.a[���3�mG�qA����\# zh�D�Bs�Xg�1�:x���'�]6'��ؾ�O�C0�:b-?{Ƌ�vvx��*�S��O���Ԩ�.�ʺ��_�F��0�l�%f��R�n�XX�v�o ��q��Gkǿ/zߎv�H�%e";�	�\5+6��!k(p�j�^�j��KF&X=Z��h����L1ͻ����\��@���h$¦S�I\���Xҷ�1��?c�Bg��&���j��w�@�Ϋ��a�͞�3:\k��󍢅m��X��6{OB��`��Kl���`���k�W�r���5Ju���B�z�	�?iV�"��"�i�T�7U{q���~��ۦ���h��A2��g�u�v��)�w,�l��9�Ϻ���7y^)�������ƺE��;�;$_�=���<-�`�.o`��k|�:?��s��"�h�A���j �|j�Vr�Џ����;p[&Ŧ8��*X��c{郰T�fb8�5@�;�+N-M��7e���Ռ^����ǲ��T�#�����<�4��|�Ta�n��Ŝ�s|��l.��Ԑs!>_si��36��qY�_�6>7�ѱ�d��Xl�͈���;6L�
7�_�AD|d��ʱ��%_�1b��e��Վ�{�cD�,�'ŪQ�|�g���.�{�ZI���d�eIj��A��E�����35�4�+����a��[[HZ[�g�A2�> ���o<�*;;�w4b�C�5�xd�f����,���s�ֻ	���6`��m'O�e"̒e��$0���5��SV �o������hn�j(��Zfٌ�(M��.�~h�D�ѳw߷ P�I���Ċ���}''�@M�t��� 0FF��oU�uu,l� U`�WHC*]�IT���MH5�{/�u�BM�g��8���_�|�����;(&��Nn����-��M�ĳ�]���@qpy��D���.�[]���׎QxKUߕ���s��E�T��t���p�@�3@ze�v��X�O�˛�j�ۺ�[����=���}���;�_�&Zvc�Wx��}�\�[�@==�c��TR:�jf�rZty��³�X�r��p46(I v10�b��K���1abi�����3����Aj�Մ,/�b��XޱRW�+��e2�K\|���e�_�u������d�*�$ގ�P��ď�-�,,��i �/��-4�"L��V��+'�U��B�oxS�w����S���u������0���O_Z�%̓��8T�9[�􃺢�0�S5?�/9���T�M�V� �q�B��햙�:�������5*4�}Nmh�2�=��̐K�q�-��9�&����{���m��@��'ĵ��EmQ�c���k�s�-Mzl��y����,H�VP.���r�E���� C.0ҰC��0rE�w6�����s�x�nY-����}����
���e2��@����~zu
����|S_QS�Ɯ�}v� �����ȁ�K-eYn�ؚ ���a�M/��Ըi�w����R  �'��K�=)&'����_��Á��A����V��&g/�^7�$}ȍ�j���;ѭa�{�)�S1QQN?����^���� e�$����||j�a-�1��K�v�i7E�k\'<:�#�p!vI�}�ؙa[N����:��
��8P�;�,�b.�QIi�Œ~2�5Zu���lq+V��3��:�#O=yg=�<W���Fsz16+n�n �3���6SR�iw����`\�	�6a41��Jfffy^#W*7��[t9�|H�UH�~����9vc�<�/U!Ä��C��N������A{/ڄ��/��D+|�gdG�ٗ����5e㪮��b��	,�j<m;���b���_�(�\%���du1hŗ $�?�:�GC��Ś���k��f���:)s�*WxU�9!�h|�~�7�Z��>��sm��PQ�S�W�]�a�d0����K:���I���c�vL�JA�ۮà{]sGĢzi:ۯ���;��� 8T�W�:����4����ˏY��.�g�K��U��r�ZA� xI(J`��%�˿�/�����qd�
��5�k�"}�_n�6*<��>�`S����	��]N�:+Nц��j�����U�(����*3��h�����QHF�p�c����]�E�0@�D�6��v��P
UnD2�ǁQ����{�l�03��-kZ}!l�wޣ
�3��0S��2���/株��01��v�������4�`ii���N��v��sv�}���
���
������bP1�)�3!ԗ_Ѓ�U�@Y�ʛ�D�S���ن���?��S�����y%'����� �ؗ�8ox�NtnJ&l�AF�0~��*�r�b���� id�ݍ������l	U�D��) ��F�Ot����&HsaEG`����,ֺ�,L�/�� �Ǫ&|���\�=FW7�x ��o��} Z�{	Dz����SF�H�����/���Մ!G;��ϟmW�ʆ{�+{�Q�	 �o+��Jy+F_�׮�c���J�mەd�ۍ�
������O�N�������G>�ؐ���7�j`���&j �! KPW���Y|d���٨x�����$a;`<|�/�e-�� ���ы��>.R��~L���/^��j*p��	t�!�6�َ�Z���] ���C\�R���ҎG>�?�@�1	�TYu���jX���d(tf���"�K(�ّ�Ӵ.�>�8+��"X�N�&F��V��7�����FqWɢ����ߝ��:��~Z�8�KZ�����uʬuKȜ@#y����,ވ����lթ�6WT!�嗮#��G)�}�q`/'�`���b�YE��xGU�B���H��3��[A����I��,�_gB����it�m�U�z?�� đV�\4����|l@6_	Od"�_Z��b��5����s��'W�=ի2P���]�3�/r��j������׋�h��Osv`�zXw�ؖ7r.� T�������BL�.m����hv�h���ߍ���HJ���I��,Sӗ!��eQ�D��wDض-5��n��Q��Y�\�{���Ec[�ÏL���n���f!�/��Q�	F�[/�����0=2���`]�3��_��c�bP�a�E��u3��V��"�:��$_���|�����S%x�j:ō�g�h��nmK�l{Ǣ�������GrL��'J 	�C�(���Y<N}�af����+�b�c�C�J�G����m痍��n���=Hd�ho�D���	J�ve���S�х��ڤN�*�MAl�Nu��h��=�$ �u���*�Yf���y&IKt�VZ���Z��KDHћ���R���ă�y��Io� �}��zI���7o��1�'V���Su�I<�Ӏ,�LwN��z����o+�^��j�o<�y��d�+֮Z�c6؎���Q�}ؕ	����9�9%!H��W*o�F��=[Vb�`ނ�b.��tU�����9��vN�Z�c���^$�o45֢�>w�b�K�����\��j�\&�m���PSJ|��>��8f���74l���҃�!��Z��«5c�|���������2�lYd�ε���ot\F�8�����3f+���kM�f�������N�6UD?��#|��d�:,�xz� r�ݦo��ʬ$�-?1^I�����E	),��8�X,��5��I����a����"��3?!�V���0k��ノ��������z���)�o[W1���.^��m����H'�bF$ot*n���L�K�$��x�ȭ�(�x�Q�����B,�"T����w�:"P�PK���J�R�הZ[�@1�ܼ� &~��Nm�o��R��[�3�(����TĦ��Ph��C���۪|��E�	a�f� m.��� ρ|c.�v�9K�S<0�XH1���B����\�%N�����ޭ�ݰ�c~��Ʌ�Y�-d���U�,)bk9�F͇�nES�D���L_`��MYV��������Y���r�n"�s�v��Q{��7W��T���ێ2�-�I�Q؛t��.���#!t�-�B�3y�;��aQ�7g	�g�6݀�՚�����&-q1�����V�HKzZU��)̆~����GEб�Ww��~�ƹ�]
�	}x��-�ly}R��я�MGS@�7z�G5B��>ڂ�[*+�ŬO,�6)з���A������w���d��������Lom�x�W3���$_�P/�nyѾ�-�Wxu���ں�$(�d5z�o�S�▆������wz���Ǩc��v#����S�	H��� �[��&XR��"���\=�V���-��N����ݓBwr vU��0H�)޷�}�#���O�?2�W�^%vXK���'�u�s4�2����Ϟd:O/s)AO�{b�$Է���Ej`�Lh�����O����z$�HYZ~��B|�i��?7�sf�;렜����iN�]��u~j�u�A�]��f�s���z�Ӻ���T��aO__��?�h�ÎsF�ݤA��2Q���L���������r%�����S6���>S`��ȍ�c�&���G���1۰[��lگ7�����ˑP��aU�p���{��N�k���c�ڤ~��O�������<�69(0�����j�"W���Un�/��i7.���0��i�f�o���?h�)@RX�r��nf���o�W��� �^������d{Y�.#"\7��c�����[z7�g��C;c,��<��=�?d����"���}�8�!]�~�+6鹎tr_Q�M���y��]Xz��Z@S�
��Ǧ�Xz�?"�ǰ>-F� ����ײ��"�2�`ۥ�}��q�QJ�ǟ����(�ӄ���1l�׈H����%�����W�jcga�B�zn^^I�ݮ6ܩzO�<�y~�1Θ=���I�~�#��ǉ\i^�>�+H���Ҏ�'>�{v	�&mVw7l߲�+�yt��x�5�TB ���#s��VGF�n-�:�1���)7Y���{O�P��>,,�?v3PF~��y�v�q9;�
����H�����z��!q�'��ɷZ����kτ����pV܈BŠ�ϵ�tK�ڞ*⠚�%��!���?���6MG�n[��`$�b�`���&N��܍/��iu�\�cF����W�����&��a������z =��5�_Z���43�֏��䢎�=�HJf�D,���ׯ�k[�j�v�;%�r��-Y�jA@�,iZ���8�����>n e��9�z=�aN�����u��B���Ri=��d������f.f�ݏ��.9�&� 2�Ҥ���M�K���ESE��‍�x���rO롚� �t�ߜ���c�k_���wJ���@S��I�iii�mSjE�ǯhn<���!�R�W�1Y�ܧp�Wc?�z8%0H�]���-�'Fk���R�DV%��� [�'��<��}n���E��턗S��V�66�V�X�=�5�y^�_����4�?�jl���>5s<X����Z˳�u�Z鿔�~�}�R�#���;"ECX"���u5��겚E�s+.L=iL�
�u�\r0� �dW�גם���x�(�y���R�n�Q�wA�-����kJuI=�z M-�����k��MlD�nͫu�{����QDF�Mq��'L�WX��jIb�Q���fKDU�4���llɡ�퀹 H�s������Ǡ���ߠ$��B2�"x�>㳓UWV^o�2} ��@�������&��eU),��9ˀ���������.��YX��,[�b�W�ͱ ;���@�|����!c*Ȗ��0��c�k��x�Ё��x{�۩<\����S�����2XX���������ǭ�?����q�d�����3�o�0s��s��-�73>���S5�g��j�h��7��������B�7��W�Qc��nݬ ���y<d������� +�K��i�\�V�4��[d�U���Rk���/{fZ�]-��Ƅ�.嘤�zg4b�CR����U+~��Pb���Z�A ��,�`l��m����E��{���t0x���QF��I�T�.������� B��m�D ��58��;��i��"��]J���qt�ĐSԎA�]W0z�{y\|o<�c��\�pPt	j��6�]��������z�,�ǻJ����yKwww5^��\�<e��rn��l3�Q	3�����}�>��i����ܒ�AL�Ǐ��rsU��_Ѭ��^>�sSXq�z��1?R�Yh���[�0��I&N��A�v�Kn�M���rzz�����	�����js�Q��Z����a$�mm�C�8�x�"�3X��ٕ��� 
�P��q*�I6�QSSCq�X���~땤�>GHG�J������ �V�����^�
���ch\$5G���뒝
��y�g��[�}q�䋛�f�@�Í�@�h��X�4*�+��+,*:���q��@�j:f����1}4�/���[���|�U�*��X����~���0�[�؜%����j�t��KU.s{U�^�%I{��f�T��w{��7m����la�4��ö����w���+1�p����>d��:ImÌ��5�}�Yq�a��^�O����_�z�;��=�x���+R迵�iqċlc��������Ԍu���#jK7_T'}Z!'�.|��+�J!�7�$�r��䤥��$�%�-k���( 	���d���V�5%��f?⬄�:���G'�D/o�5�_8�x�r��4ܱ�����eK�^�v���y��33�:�T�?5��{,1/�ޓ�U	�Y�����Z;
��3�����E���-!%%®���Pm��Vg��B������I�½���s��q��^Ï^���H.���P����o��g�Gp�q		!����ʳ��E���� �⎉IXII�3J�4�ђ.v�k��қ��d��(�rK�_2ه��o��*Q�Sl�0x�����i���$�R�DZ�U�V���RE�{�+��V�Z��v>���l������ܭ5�`�3B�q,�z�w �,�Ҋ}�7��L���OB������75�pD]-�y����?��a-�MB����\�g�m�4�gI���n4�*����=���ZZZ.(*�uvvfe�ɷ��ի�Y0�J�s�����u�oM9eT���f���-�����a�{$y�Y��L�:�1�o�%�Ւ�Xl˦��[��Z�́y���/G#?Ǵ���ې>�k����#�$�g20������Y��O]���a�
'�2�w�^x(��S+�������Q+Q���,�|Z�d������8pk�L�s뻓&4Nf+�9�}A���E��*�8��"j���ot3c�8��r���%U���e��Q�U�Q�JSMr��8�{��e킄�QoB+mϞC|v���32�Ԑ��O�d�����2�6L4Ѽ�ƻ�ok�~֑�#��'���߰��7��WHZ�c\+�4��|,ޤ�,� &eڇ���ҚӶ-1ȱ,����|�ԭn�y�dV���7��1+JAOO���]����<OʊJ��Ɩ��Չ�y���z6#�����sc��n�q�7u�ͦ���+É�p�+x恻~~�D����A� !�+�: �w��w���&.��M��,�<{� N ��˗/�զZpZ-��oa�˷�S��skAc8���U8#��~1
���.q��%'�C�K�og_;4,|kq29��=����rs�M��3�R�<?/�fh�s��l�c[ˣ:$
����@���>��"bb� s�r��Wa���/�)����!CE2w�0HU�@^haOv���Q�����-�Av�¬&-+n�K8;:_�����NEܻwO�={6��N%y2˖��i�C~a�s,ek�v�.W��
�Y��ab����W�6��3�r���T磤6b�C$�}�&a�G�x�}���!�ys���h+�$��Q��bά���j~�Q���f^H-��. I޽{�q}���a�K\ ��j����w��o:�M)����C�a����_��	�T#�b�%䖏�}1�=Ck"�=/���������bG����3Jv[^�3�zb'��o߾��G;*D��85��#��&'�4����0�g�<�u�v�����+,,R��4Ѿ��vN�F�pt���`��O bW�����Qa`@����rc�4�8ʅ����
 ���Ĩh��ZP@��NV�f�m,���퉩�ߪź���G���^#��/�ﺪ�g�t �ou	�� �\���E�:��f�x21�7Pbh9��7������+[H��z��n���gj���u��n�������W�C��FoAQ0�aÐ�k�SnhÐ���la�QHH�}�8c��P����ʞ����N���8�AMQ��S��z�W-��x}��.���ﴚ8��}������������Z$A��xǻ���a�d�Բ-�/�R�e~�>��X�5�]���A2S7X�������E,>�aq�-+LB<�=����侒҆��������6��F�9��) Yl�N��d>X�هr����:/<�BO�Z᪜���/Y�E�D���� �jQ� �x�&v�B��ꞞPc��I�:���}�T+ܭ�L��3����<p0)���55Νw8�� �+ck���j**�@t� R������,GH� �}� � T8_���]轠����"�����%C4�da�{0z�m�q,���aPJS5�e���v%�gW�ΦzaU7���A%���3۱��&#�/�J]T�P`Ϫ���X@����I�3�?h�J���3�d��ƈ�rť=��i�Xa�`j�2Ȧ ��`P�T>���'c��KROT���!����)~�$nhh����QF�<=���5���'�{������RG���qVV֔�,Tg߽����܇'L�����>eq�߆?��%70�w\�e�~)έ>9���N����R����iQ^6I����qhC��k����(��F��z��Y:9fۚ����l�݂F��q����<LLL��ߟvc�ݵ˳Q���N2l��[a�߳&i�?�OOO�+�p|NNN��o���"�CG���'����j��
L�6�m��EDE�+S�"-�@T#k�
�9��WD��&���5���߹� (̐��U^���8d Y�	�sf�>e���P��6+��TOl����`�.OUS�����?�Rj5q�@ � ��i~,����a��7��1��<iI�:�z�)��⒒n!�hT�·}�u��_�ߚZ�s`8�����E"@ �K�o�Be��گG����YQ��2�0y�jZ�Y2���G �D��d��T��k���֗5<�$h�#�{+k�qP�X�E<�Zl���a�XWGV��i��	o^����������v|��{=�H[uY豧A]:��w�ʦ�j�Y*��O�t�{�?�����9╈8�H�|D���=X�7/��� ��֯�� ��[��� �_C���w����A���B�u�ss_����n������Dm��]�[�ћ�4ջ�z�I��^�4�V�i��?�����u�cW�Ɩj��8;;�o� !Y8v�iz�ˀJmF�����ix��)��ut�uA]�\k�0_�&k���n5z|7�#�ڇb���w�xc_��%�\�R�o(.^�|�q]�5�$�6�;Ge}����y\T�n.{~:�Ԗ?_:��[<rDZ,���Ae	?0x�%�(�zV3E�GCC#�=<�ǁ�����# *1��f���6�\��tFJ�J�TMaZDs0ϗ��!þS�qI�Ͻ-��]g���-�f�f�h���>�?����|�j���Q����U�z�ɓ']��~�t5#��� �,�<��(�}1�O����;���<��7��Ж�OD�ߥ}8N���Ji���xd#GKj�������_���o��$�Z������'즁 �vu��J\N�8T9�����G^"Tk�[�kc����uR(�C9���eCG=&�g8-��%S��g�\_�ʂV���X&�4�>"�X�٘ά�?mm�|�)R�s�u8�X�^)]�Z����:�wC?眪��|���sȩT�SҞ��=?�Z\���<������Mc4�d2juZ�����S�����NP͜�q�RB��g�8�g-u�1#�^����\�Cc~���'2�(�[bh�����P#R�$�i���P��^�[�tV7�j82���I� �˪R�6HƋAeFf����?�mIþxB�R��IUO`� ������^�Ǉ��N�҂ZG���E���{����;�f�������^�H�G�'�������tɆY�ʛ.6ǂ�M�{k������+..v^�9ruVFӸ7/�r-�(t�W{2�imҸ#��q>�΃Y��U���ￇ��ݦ���dmi>��Q�]�h�@��l)�����5ӄ?���v�EMǎ�9�Z�͹��<� �Z����i���i�ֳi����'���ܠ�Qs%�à���=f��qy�|�$Pf��O,sYJ�����|v�O�����y��S���o�/e��OqWk�y8�0�mc���.�zs&���*�-
}H�p� -�ѣ�O����v5��W�J�{�=҃�q�y���pImw1� ���x3z2�'U�S�:Y�����/�kci|����Ȭhe��E��J�4m2+������v��tܶ�����R�Ԅ[�H#*�˼�q9lx9,.>��PwZ��U�_�&�r|�[�-�ٽ�0C;�n���иAGW��@��l��,D����]�'A�0c�㠼o��l6�[V��2�K�	v%\�x���Γ_����7�u�kY)�Y��69����#��1�ԧd�"B��"R�C�Mm���(5��b����*	���e$_|yV@@G���A���M�ɿ�k���}�4����~˖T�	]+� ���F��p*e�V�	Y.�R6�R��cKT��b,�Ĺ d	5�M��ZB��C���o����dC}+i -%k���l��j1�j�Xn=@�윗mH	uB-&@�aP���P
'LT�/���x���C���:@}pG�B~�P�L��d��6ķ.����j����u0aF��L�:7:\��7p�n.�D@��Č���զ���,g�M�w{4ÁW� uP;���e�xc�s��,��kk c�
�D).�R<"!!a�L����
��>#$f���/C��\��@u7�_Wv%��]�{�Z9>���C��t���tu�U$U,��t)c��~�>ǒ6Lt�����$���<k:Z,��YfNR�S�xz�1�u���I��9��M���(~"��t8\��}]��H7�u���9�^�A������r}�Qk���V�j��ҵk�5r��lWb�d������Ě��q@|��Y�����>\�f��'�(]��C�uکsp�
��dd��{�����*�G��D��������Llu�G�ŧ�R�_/n�(6о�Z�y��XXǴۭv����jP���ɞ{�F�+k+��{�Ng��6~R��@?��y�9�幊���ힸ�x���?_���Ԡ���
�L}���zs�z3��#a@���A��VIN֍/ʦ�s�T��-s2	�K�飣���4�S���w�� �`�����P)���&��;�1� 8@{��b��HD0Q�I���&6�E(T���{�Q�r	5�"3�o��������@;��t�����O�BV�ʹz��'���gW�7�T�r�,�$=��fiZ*��\��&M,�<�s��L_ĩ��V���r̷����O"wS$l�:��r����$�K,t�?�s��U)�Ǧ�Z�|zu4�v(0�@����Y���;�eW�4����9B�<������zM_Z,���ϧ���jJ�x]`$S�ql���1����-9(�%�LVg�����}?�23%o���Z����1����I��C��NS��=��-�
��s�y&���Jg��5�PNw0(h�t"?/ʃ@R$����5��Pf��!ⳃ{�X:Y.��� �ۥ��#|J$����O��X~�M�����:��qZG/�����6�.��d�������i2���nK�+;})����9�=�WF�m���hW�*n�$�w7��X�KY��֔K�K�nŮz��|�.u������l�ண��`�B����$��R;ڶA�� z��|[i���&�Q�{���&�)_X�# kF�a.�jI���XW��j{]ɝg�C8Vb7YdF�,�1����@P�F� ��vhVp�8\��-�k���#aW��8(�����q�n�X�IQ��A��V�H�Eq������ZN��'r_i�~؉c 7�6K���T�*i��p{{��l�0+}G����Vּݟ��� ���~cf��,J��ł�`�	�9�Q<L/�ޣ�(�	�ϟuwQ��$h@�=���l�V��s��z�P��r��|��������� -���
H'j^����j��>����k�8 �ɩ��/
w�K�%D��~u����0K-���F�{���gfz�������V���zO�;N�y�ː��n���(SS>�F�E?�[�H�����w���4�aM�y4ǁ�g�s��C�$����,mcvBLE^c <�JΣ��|k�i]6��a���д����u��2������{!�uq��>¿��!7�
��e�d��V� C/����$�"��7�g5�@�ǣLC����&t�zz-��}B�	������q6��a�|�E�E�_(w�5O��5}`�7.\�8�����$.Q��������OǪm��H����b���9�$s���ˆ���J��}���u����&G�E���޹}�������|���X X~}qx�e�Pf{��w9�
N7�!E��&��Z2�0��2i��j�}�"-��t�Z)��IF�������p�8��͉��8�U�9��<�1H�w����7�@iY9�k�Y`:�;ooR|}�C"p��������{��_�p�ۇ�:�9L�R{�)�'Ĳ)��sM���#Lf�Ч������0�M:��:�3c�����SV��ؼQ~�#?*CB(U�p�qߓ
�Z`�Q6Q�?�G�.�|�b�}h�ҜҼ(?�6D��W���`�r����b4t$e�+c�o߷5F�@�^��Xz?�>_�Yo�pgh&��4�'&���7��V*�QD
JY=T��{�5�� {�:?<�qV���l`���(>@$�Q)�V_�|�������X�T���elvP���/t����:UJ��pEɹ��u��������d2��{L*����Y�#"P?�.��I�C��_{YN�����[����9�&����㧠}U���o � ����POw�*n��0��4#˭��GmN�+�ph�h�aL���Ŷ�U[ĈJb@�X���a�C�?@�u����M�3�nt=�#�����#U��(��P�Ba���[N��Ү	��ܾ������R�S��n�4�M��k�Kǫ�o8KU�̲5�"�C]*@�$�g Ԫ��4=�'�"�^w�<�R��gT�C�=Xr^�񰁲G����@����t �钐��\#F�R����Hx�����XT.�������<̬�1�^�/Ԡ�!������5!}����T�>�@�����;*����G��/�%���PC�l��-~C6�ӂ���n6�4���h&��,c��{�U��>d����),-��0T�����nV����:����8` ���J+!ҍ�t(J����7b R���"�ҝ��|4�9G�}�13:�{��g����}	Wv�J�Ϲ���+G�r����Ε�z����9�[L,�:�]z7ތ���x`�(MZ�h9���(8�!�e�(Uړ�}����W��Y�̜ӷ�5�cF�CG��_�Ǧ�al��~���<_�ƌ��m�
���L�kf�z�<
%U��5����33d)|����"��2�e֓.��鋺�|4H.�7�t!Ρ}�I~�TSڇi����˼3s  ײ��*}E)wo���<��&L�	���+sg�=�����E���.G��.����@�C����>|����L���AQ�ڿ���ڽ�t������t����1
��0@2����i|.��T(�LޅM��p�'��*T���Xl�8_-z����:D�Ft�\�z!�yG3��q�c��˚���鎌6'���Ά��4G��^[=].�bJEW���ܟ�3�d�`����:Z��u���^@7��a��h�V
���s���̫I4O��B�++k�zEĉA����q�g%O�R��q-7��_J��S�o�#�P.~�"�t�i������F�ӛ�&����s�[�pI�>r���g0�x�
1�y"��%F�K���{������VY������2B�\���~Y(�X���>����W�����3��3(HI�+*�iJ�[bF�y�����J�=�n. c���<�����`��ݜ(�j&��YP�9�Uq�=�yDC�/cu�����-�g����]O4��'�_��q���@�a��?���xj�9qJP�i��$������E2x�#����?�B��H�n��@��i�&��8�'�?)c�b����{���q-�P�FѪr�����g7�QJH�}��D!�d���Ν`�`I�5�G��S���(-՛�<�U�����o�[�ń?���w�v��U��+�8�9%�}�{�Θ�/���|5���'t����s���[�C�Vo���#==��=��E��/'�_���@{����Ϲ�O��%EP�44
���S�^�P����X\!�"���}�S��?Z�o�X�/��j���	�qs*֐���U��
`�?�f(c
�ӧC��8{X����p��L�	ǿݟح�?4]7l��$?��%�8=�&9�Ԙ������Z�I�Ac7'�c����w���{�A7"����Dߠ���� �*1�$�# �{�6�O�
)A�s�ǘ��F�!��o��Kmd�{���g�p$F���^��"�����T��+��Uǈ�X�O.w<��o�Fy��,�W�(B׍���mll��A]|'<m��w��P���Ǐ
�I~�eW�R��ZXK���w���$��|���ǯ�X<0r�����h�ې�#�F4G���ʥ1����k �#1��q;?W�I��?mF��H�����vPZV������叼���K�����8$.�LMM�_��^�3'~]�.X���㩮���K���iD������S�.��1 t�Ä����x�?�(�_�O4|r	��,/yb��`l 2�W�
�g&��E�g�_�H����_�;X1�b m�Տ��~b��0)ݥ�/���L�)�$�	����'�[NB�ĔB�����,[t)f���C2L@��4p1B�<x�_�����w3��S��vs���IT{�[ۻ9}���g>������s񧶫wmd󢪼������h|��A*�}
Q��XUtH*�K�Li����ܿN��K�v9�b�zW�"��^�g��{Ebl�,�Ѷ�[p�����h{���Ύ=�?�C6� �k�`��)�B�3��X�}��������7���w��%���c�|�����:�_�׎MQ긏��5��7g�h����*��}��>�^�3���H�h��-�S�d��"���X��LT����D! ��E#�dʛ?�T�[i�Y�rE؞��Nl���ݪ��^��|f��k�	gs�U#ມ���Q{Os*��mg�NJ�_!a�A䤥?M��= ��qΣ5�z�bh�?��>M-�U
������������\=�@m�(���mQ�����`dP%��~|"jƊ;��V���<+�yo_Q�l�����F���Q����.����s|���e�r�	o���n?������'8�
�=�q^ws�.)y�S��O���Y�p�1I�*X��@�������ޞ%V4~Ś6ڤ�rY|2�5PK{z�Zm,��!�w�����:�9e6�<�.'�ٳ���W�:=4K����Q1���%K[�AE���0A��z�,��)��+��j˥��hnUUU7n��˥)RN�aS=r�p#?r:�d�
������ně��ρ�LLL�8���������dq�[�U��x3ʈ��ܨ[��|��iT('p:��mjc�_i��{�V��U�:��pǶ�WL���򮯔Ebl	~�c�W��L����".O|����aC�3C��I�yR��;�_�ʲhr��k5�iB(4�6�������I��g~�����ʂ�1��S���7���ta��t�X�q)|ic��n�=���Fd��Բ
#��݋��*�)�L��7�^Bң���cD�w��L�"o j�*��bF���t��Ͼ{�̿ŕ=.pl�a�Xm�i0���XNt���{0���|~ �7�j�	T XB�g��4��a��(ț=^�<>rx�ݰeP�?�����.�����N�J��
�ɝ�X�J5@a�w1�b�ZI�O�{����}QJ��������'�$���f�N�B�Np���������9���-�c�Zr �l�y�ZG�E$����eZ�tdCD:W����-v�!k?t�jWFJ��葹��L�C��$�ɽ,#ls0-l<FH׀�N{W�@V���:�2]�{m���
9��]�v_l��NU__�(ie,�����20v�]>�K�O���o�?�g�`�,�waa��z߮AtX��>�{.[[Z�[Y�����w|���%�>8�F2Q!~K�6=V�˭�W,��Q������:���:�^T����NN����4�!�O2IXGI�u��k���]^�
Z}#���R�VG��R��d�f��Hd��"�o[��0��#/%��P��y�_�մ��h��}��h��w�R"��N�����e��S$l|��Ϟ4�k�bh���\��M��o3 �B�Ώ�(;�C��-Hi;[FY�ݴV��~����h�y�I4:�")!���B�&x�ɀ]d�(�Ӳȏ��k�9���h���Yɕ���^�K�Ofɳp�S�#�#��7v��;a$�T�q!q-��H�~Z�@	�W�U.o���,,��:�����=D���W������v���\���sєm X4ە�o�����ٹ鿊�� i �PY�����3�+/N'���t�j��J�	{���2��#" Q�~�����kR�Z��Ĝ���H"�H�U��]T�{�=����%���A�5��m��#��&��犯�� u��׀e#��~�I W��G�DA,�>�}2�����)?��%�3�om���npӚ�S��z�/�҂Q��P���.�󈈕o=O��FlĴ��)))����>�_�FI�(��)�&v�<�qɛ�[ct�wR�*M��_8>{�JM����|g��X�Y[a@i�W~���*I�r�k��el�>�Ks�+܊u�q,�d������"�V�ڤ^�'U6���#�D&~���৤�v�������DI��-VF���1�� tH�9��m6%��D�6�|��KA����+�,�İ���[R%���N�g=�>�O���T�PQ�3��!�)���b_�bRXU�v�r,��e+��^��h�PR�ET]YO*�!�w.r|��E1�#|�s��}�;���K1t"淬���R8o����9��d���ꧧ�א&�jpSiX�x"���n+�(�	ʫ��s���8�#����v&�t���#a�8:�x�%�<��<�R�1���ߌ��c�[���0��\��ؑ$�����R��� J��)�˲S|���A�ޤ}S)�)lon{x�e�\�=(C��S�9HĪX�A����w�L%ߤ��iܺ��l2�S�Zl�d��Y�1_8�Q�:�0�\���\	H ��f��� ��oVa�U��k����5`Mϙ����gi״��@^����1������q����p8U�^3V�7��|:;;o����3�By�~��{�����o޼a��!���M�6+9l}9�w�ŷ�H�"�Q���få-�tzS�e���:���0hw��D���	\?S��'Ί�'t5{[����6�nY^F�5p?��%2�&��T<;��z�D����RRo�H��?_���i�j��Jã����DF��xFr}�v{��~&T�0*�g/j�;���<\'A�V�e6�(|���S���6�����#i2,�F��Q<��ʿ�X�i88a���׀���
b�i������?����o߄.]�D5���<�|�aޚ�Z��=T���0��Mt��ė��_4�p����D�����&`�45���?�d���XU�	|OOO��(5�V�܏�������O(عקN�E�W9�V
(�4��ML�
���+����r|;m0<���O�Q��؛�;��Y"Q�pvHW/dB�`dI �Wq�S�V�94@�o�W��G�@��*`����oxXl����+,E�b`@b_�xTV	�N�1	��P��*���F��2�Zi�]���7�>�E����s�oܜ"��xԇ�f?����r���QP�6 Sz3�=cc�~�Ǣfb��?���5,,���4�4L�"������*Ww��;[�ݜ�V��,~�I���`(Jf�r12��/��x�v�Vo�M����^H�=U�P�Ѐ� �_��U���k�S+��G���$?���s���;m_xt4��.Uŏ���>>� p'7��� 8�e��	4Ng ���k�H����P�L�p$Vo?��l�������`��&Nߘ�	p����O0�b�1Kb����(I�`(�c�1������Z�Ͷ[�:���u�"2@v��,�%�������yˈ'_�%@�G�?�]�Q�!����\���E��F����i�Vg��@���"K���D+�n�xC+k�Jn�z0����y�]g��*�:@�;����֖>�I��~����4�Xy������a�(Z���[�ųE �uw�gT5�m��V�v� OO�yN�ֽ������mܝT4�˫S�Ẫ��5F$����pO�aD�X8�3�p.ΰP�z���e=Y�-�/�W/�h��0{?%9�,(����.�WE�Ҝ ���6	�K�v����Un��K���	�k�G�m�fp�a(�(V�0��2�M�g-��n#HͿ�3	��D��Ȼd`
@�8nL���]Z�"�����\'��+'tlw�a���� ���p�	����0�ӡeV��1cw�骒<�eJi���6����0���m�&�ݣ��k�R���t/��Ҫ	b�o@J�Wa֦����2.���b!��+S�����CN��ҳ�����>`�+�_�Q��7��'��PKM¶b���^ɿ65����$�U��b$P�vFن3�[aY#x�e���]��u^�d@��dɜ���rC�~�9���uK8�Ԣ�B��ۃ? >�7�.L]U�"��0Vy�dƓwKV�3�w^�m�%��%�NxCx9M�W-A���sJ�%c<�.��LG��Wp��WYۧ_	]=^-�>p�7oz� ��ng�cU�6��!~�&E�?��"��ɇ'�!w����Q=�0b6fĉ{&�y�������G��ἃ�>�آ׉)�T.�ۛ�ةÀ��ȝ�b���m����+/�2�*�`J��ư���҉10����^��T��#�溜�?�{4�;���4�|2��M4��x� �E���CL�2���� W֭)\w&0�� ν�8��O9��H��YXY��*!2������� �Mv������`��ݓ�h�ĉ
�k�Ô�Q�1�?���E��VI�,��������y���W8����2��k�M�l4,��Zx�e�w�C���es1NLG�����o�H�d'�b���
?]����S���.�;6�s ���i%*x"7̏dZZZ�O��DC�!u<L�,mÉ)����\\X�-$Ϫ<r�j?�F��ϣ�(2��DH\\��8�E3p����J��WC}9��CD�5"dg����O�������lBu���1��X�%�u�e�8�ʪ��y��vF���ʃ k����U��KFڌ)��K�ٴ���r�O�s'ФK���U����Q϶�p�g><<�p�Yu��<��O(��sh��	Ɏ/x�9�RѸ��krWýV��xyOV
nݓ�F�c��0�	Z���gFd H?�,5,�H1��چf�]�߉�ӽ�����FNL0(�YM��'�L�=F^T�;����ɨh��uN�K���h 3A!���e��)�4S�������)���/��%�$W�~av�u����xYu_����R�����vK	���'�Y�Ɵ�0��j�fU�F����tX�IJJR�;Y�R���V�IOS-G� H}��#�~}�0]57I������0ky��F~kkkA]-��
e�n�Q'��Y�y	���^�B{0M��� ����pvو}�᧱�D�T-̃�!�������f�_#�Oh�����(&Y��
�7p����z��������f��ҨG��!����
��ȡ<w΂M�Z�X�}Ç�Pz��HX�Dg��;���())Y�������T� @�@�-���)��� *����͘���)|��-ǧw�oPP �W��f�@H@�|����9��Zul>���I0��P�0iC	Gp8�k�Y@� !<cU��%U) ��s%����,,,��0�঩�j������<�W*�0h�GT���߹��Yu��m�T�,&ֲlS�~������մB�cxSvvۃ)s�#�����R�<S(��K?���Wa�--���ehs�Br,9�o�w�꾿���?�Y�y���XPR]�"���]QQ1e����w��q�>�������OᲚ'�wd�%�%��K�����_y���͹rIDk��0Ze��C�6��x�j��Hf�<�?p?�I䱻� ���/��u3�ݙ���^�J��!���iJ�۸i�25nJ�2� �G=i{�^�	!��zЄ�m�``?*�HR.�[Z��3�V��D���Nh;�	Ǚ�`˕⹺[��H�m�Io��l�9{6)�j��ȣ�<܂;>�F�yc�V��v�t���F��_�<K�#��Y��ȴ/]bs�ohL�gȀ���(�.[����35�f.��������!$	�PFn�{:�̻���isb�3���{�7��Z�"�S�N
�����V�py�_{uV��~g���Q��"!� S���8��~��s��e�M�ਊ���i��U�~��R�G;�h#<�x�ɽ�29�[>��-��� ��nh=���_R���!���	�!: y�~��0.�eve�B�u/Ӹ�9`f3̆v2��;p��O~�oyGu3�?�(�=.ג�D�� Ϋ*�~�������VF~k8k�y�ȝ굱�}�j���$��fpMܴq�dr/��9^ '0J�}FG��2�j�	���e
)5@d���-���\���]�?���u|����ˀ�T����LWɾ���byp�!\ R�]�.�[��{����d��O�za�`�)�=�2E�P^���x/&��5��gr�i��#�I��؆�������aY)))��K�d(�[L��if2M�(�G��z��R�z���<���$��[�l��%����Z/���l oT����8C��c�^�H�嫵��;���T�n���x�4�G�hJ�mzI+ĺJ�KU��J����+�*vΣi���ǔY���ˆ��ٗ�y���ck0�ҳ�IGf_�/%�,���hڔ}����?����D q��!���X2/"�6�:�˗.�<Sּ�%��8jhkk�-�.0#��s*+9cL�,AL����R��N jw �:���|��oŤ ��� у�%�}�� �niٿv��^��8�����5m��A�s���0p���Fq��;ڦk��o��@�M�=��T@�s}CR��A`�T��XyU����Ƚ��01U��7O��zS΋���u��?�Hk���\��D���� N��W/�ڢך+�ã�u�}w�+����>߮�%�3b��;ޔ�l|�`��=���R�`sӬr�����
�C�� �ϩ����x�4}+Wf�������gv�ni�0�&᎟Wm��'y��j��y٢��1�� H������#{ї	�y�VXJ9V�҆�5/
�G¡�W^�+E�p�N_a�u沟�}���`���))<����3#�c�)b�*����	hJ,Lz1�BY]4=�� ������1�����Bx��i{%
@�s��z���Ay%ͳ��耒!��4��[�+��[ևʶ���Rװ��;}JH��s������o,��
�<on_9O�iֲ)�+�ؔ���< .���I8�&�PY楫d��A��Yt'w�
�U�1���ܲ�˸����Z7�cH$�����$Akț�҈���P�O�K��4鳹ڽq�8.;'��?�/lߪ�g�<N׮�[��/iVBoV�@S(����Ė�������(�򞝶?���8�����!�-�?��=Z�MThdk�E���#���g��?�"��:hʪB��~~���_m�����K�5d^Y���Y��(c�B��<�ǵes$/Jܺ���HY��ٰ������<��w�+�`��fn̢�2ΊLSw�j9z�gEY�A���xO��k�,YL�F�9��� �Ɠ��.<�Zkۯ�0����l����ape���ͩk�\P�fCL����E"&ov�>=2]��	��������XmF�h가���)��T����ʅ�M��Z�����Y��*f�?�VW.)�/���&���W?��>��<��NO�潸r���5H.��|�m��2!�i�i%a���F��s'����l��u=��+��}��+x��0�x_�&ȟ#&66lf#����s�w�T쏬�u&��6�pq��װ��1D�����W^���m%���P��!Hax�RN����~�S��)�b��Uܸ�Q��0�f"��+7�@
�q�vC6A�ٿ��hּ���>K���Ę�yQ1� ��7vwJ���:��Ƿ���4v��)g�B�T�1*`t�/D�2�t���>a �[��E�h��sb������G��7϶FN!�h�PI�m�y��գ��:��.f��Y��������@��(��/9u{x 	y�s6�#�ݒ�h�{��g�����+x� ,� Atm ���i^��1����նaw|���L:}�W"94r�Jy��	����w·3�&?��vԾww���>Ё�N���h�>7UGb�_��o}Cp�S�F�s�g�:��~mr��x)6��&\vv�΍��=p�lӯ����>y���7xk��c�żnw��Mڦ>`~��/�:-\+���`v]��v�]�&V�ub��OM˄D��mU��n�aiI4=�æx؃ڒ^/}��o/ �_��h�A��	\Cǣ�h^�]n�����2!�7R����9;����H��4���T�.d_��� �R`�����l��8��B��m�z�]Cm�2�ڸ�0G�a�5���b ����k��.�Ԋ��YZd���	1�ǲ@ɺ���i�7���>C�",#��'q"78��_dn��aM	�F�G�>O�� �����HӰne����W�*4��o�GBr��l����������'� �HG��.>>��Ȫ+:(���P�.o-Z�q�%�t������Pa̝�I�;\���W�E�aְ�A6Y�!qDD�f��M2�yE��RXp�� o��$��fn_�*>������<4���e����h"Fz����������u�j�)��m� ��Cѽ���@{�M�(c��H��Ճ�հ�+�.P8��Č#⺤Dn%3O0:"�?2e�5G�9jO�9D`Zf��7�\iƩ@�ku�x-	)�.$��Nv��}�g������RˠQ����iF�ؐ�i��1^���
����������F������=�@����46�[8�E�����/�pp�����2{��*\9R�!w$n��>x]C �+%����-��OY�k"��b�X��"��ߚ
B11jB[]]W#���r��9�����A�
�:#�w�b3lv��Wc��dx7ZX�f39�_�br�Őz�G�v4��^�,��$1���0)�`�0�����x���>L�����5��� &��\�;�`P���~�D�ۓ�F<EEE'��l�Zdp4z�R�ee�7��Uz9�C�۴7��e3ca��0Hr5�u��ָl� P��m��G�0�%���	�־�ŭ���@��@`$��#��r��̤�$K�����*��Z���ȣ{Ye��Ɇ�3�n�jV0�$u���F`}sB�PR�D5���A]-c/W�7\e?�'�l�j��_��]��U��32��6~f�?��Ғ�A3(1!�)V�~�&t i��H.	���I/��c��؋��5]h=��;�D�a�����l�ƀ��B�s��>����i>R���lֳr�0���%���>��.)V�R�a`��J�6�����f����vK?�vU+�/|
�L�qʫ>ٝ^>�<ރ)8�sB~o_7K�%����#�^<�vq�#Iu҂��b��S�V+#�j,p�?�(< �͛�J�|y#�/��;��=r��oe'��Z���J�mkZ:��:��}�9jO	�ER;�_�N� �f��n�	;���w�>T��A_	�+6�mĴK��%�giJ����m�L�O�r��~va�1ypd������V���v<*	�p��<��f{7y+� j���cm�G��<[�M66��9vso�^�W���D?�`��N*�Y�{Y�C��0_�W_4�0�ܿUQQQU��<+c>V�e�󹴴�����#@M��-:�k��
�]�+78����_�0 VV�n�% AM
v|M̗�x�[Y�� E~��)��pOx`�iɩ�-��Уp!�q7�ug�e���jy6x?�d�b@�wc�Y��M&[��:iQ��se���&N������Cq<�܉q ��P�ȂY6zG��.V����!��?�˪��*�#"_��Y�H�,-X��������3���T�]x��P����L���] e�^�¯�Ў��YǭE�d�H���E�c�4�B����&6��`"]8���,����Ua��`�P�V΀9#��ŉR������I��a����Ax��t𦮮.�DN����U�v~tc��]g�9a,8 :9˞R
��)�9
^;�
t�j�5�NX 3��Q�&���1��d��Ru���'�����jb�@@&�%*�C���&h����}��_YC��1 �
��8������>֬���L�'Xsd��%و}0˶_�5A�_���B�}u���_�ឞ��ɂ>0�`�	���N�<T�<S�\I�S��3L�^t�^��d�E�CT��� p��,t��M'a�$�ŧS@U�4*,�#9��.���=��`+�J	j����˵O��T5����-�O=�����Wm�f��|��A�d��b a:�e{�G��2�Jp��

�#a�@R`�2]ϴ?�\��7��T2�P�:TȌ�S��ZԂ�#\��$g��i�S��'�e������2�NM�z�G�N�~�<��R^�tӠ�ׁ��B �}��+�1�<��do1�=�#�P���!�+��f��4�<ű�ű^�x$������/K;v`�����Z�@L�C�E�)�����	�%I����v'�$��k��⸀g��/�l1R�����+���*�zr���Hʻ���������!���� ���(z�}�Ԭ�@@@l��Z��a�g����rĶ�V�r�Wd_ê����'�0�44�'(0'�TO��h�����\��hS֖iV9�1(z���@.�j� �|�������*atΓ�����w%�1���������Ǉ@58߁_���<`m�a�&�J|щ�]��{�1"�|��(�m@�UX��w�ֳr���K�w��;�L R�(��B<Z	�e�q|a�%F�RE�'m�cb���W��jnG�ep���m�"���]�-�7s>�W����&%�>�{.Y�؂���keT�_�ɥ�=�pr�ʕ�$���6��g��Qѽ��SA�� �J'{��G��Η&'�x�^��R�Ղ�g^�ߺ��p[O(��W˴�$��U~!s~��)r$�v�n�������g�f��~�9w�F�������ѧ���e�`�-�[��c�Z�7\˝G�[�b�O���
��InOT���v�O`�����ٺ�#f��?QQ��P/�T�#t��q�\S�C�GL����?�ٮ�#�B"��'������5���4��~�ݻw�K��o9�!줦S��z�OU�V�fS����e�|_�2v�\�8.O7��m����@���~f�_����s��y*�_?&�w?3*�����$�Os Dn��(cl���Y��Ͱ��բ����m���x��+ ��6Px8/V/��%��^��%����A�[Ax��42��t0E1��>��3����v��f���ti��9��5o�{z`~�z$�䈬�����}?�VU�Ւ� ��}zZO���'�Z��}��r������e1��σfK.��N���	0��s��XI)�=+���ۛ���~w��R
��r_��
�!�$$��D���QPT|�ev���@�d�0��Er�'����b�w��4��������_��
���SZ�;����?��rr�z�o���J�c�2��P�RC���̱~�ve����K���Eq[��LOg��1�

�ҥ1kU�YvF+�$8����g�4��O�ӓ�Ѹ,�A7o�xR����}yE��mQ���$��О�;c����v�]|�ý��'��F�&�J�b�wcw���e16�"�������b�;n lc7_1Y�Yv��!�ub��ѩ��_����g�u}���/l��
I�b��b��j�Cz�=ꔚ����b�i�jbw.VLY9tI�l=������	�\����O|�^��"�z�*������^�(ѸM��Ǔ����ss��z��n���פe�=��k�����E4���e�M��r��<�;�Bq6��Hd�d0]5��Ƞ��7e�2����'�9�LG��͛7#�T2���n<3�\N׮��H��a0a�w�:D���tHk���<��岗��ewcn� a?�g|W�:eq�$(8�8g��*�K^^�CV�����g�epD:���S�u�x�`�]������N.��*�%��[�;�Z��Dw��K��Z�+�6���3G+!!����|�)��@H�������-nn�@�������9�����i�� ��p�O��d������~�;w��?I[('TE'+�i�z,����#�@�>>{{�Z��vϳ����C�� �@�����.#CVy9�y�a�W>�/9����Q��z	�ͬ��0Ad�\�Pi>X�]f��^�������9zwKMΧ@�!�Ԛ�4��}_��7��V�� 3����%�B�g�ࠠ�f��e��4�;kS��z��z��>4�[[����u�����!��ڊ��� s~y���jƪ�����À�G�}]GZ �X����&N����+Iҳ�����@ͫ�7>FG/#b�E�,z�J�H��񷓁�9\l-��HI=F�������&�S��|y�)���G�N�d-hKp2���G��`��������EN|�A!!��Dېރ�hQ*0�F�(�O�W�fS��,�Yٚ�m��E~d�JoL���k����+��.���|���	��B0r�=�q@��C����k��C�����?j�o���}�����=/-���{zp��F�zz{���ϰ��sYN��>��������Sw��Sa��l����*b6�M���?�� �/�_LS�RJ��&MݢXCa}����i_��yᐼ�B�^ɳgόLM��,��j;Qq����KI��`�#w��i	�]��TOh��~����06��Sw~��?x���D�����Cs��"��c)�i�;��bD�
���I���)_�0f���t�?����"����|��3�5.9����4cp�t$s15��Խ�L��O���m�� ��"���f�>�����%�P3�u�J�	Z�]�Q��09t���y�u{����АJ���E�}	���Z���=�ѹCȬ����X��-�Ѷh^ve;������ě�s������ױ�r�+�r��B�og�����������ք�\�����+���]�|Y\F��A `�Ց�)�X�߇��x�J+%�@~���/,��p�}-.++jo_��+�����ެ8���L߿'(�j^E<ztX� uV��ܺ����X�tv�-7_���}����	� �E��%�ύ����
G�����HX�'T�_���b29I1g�LR��
i�bj��5�GKfB��wQ�8���M�U� ����Bi� 81��{��Ř:.3S־`��5yw�MIoc���͊t��@ ��2Qo�K�#�3�P׏�$$<�.��1�� �dt���e��]ji��]�䤤�AA�)eMV�cS�G+�]���F����o�J�Ej�j^ơ��	�ABFF+ bC�و���cd����c`�YuE�rE�$^���x���8�.��o�������Çr�ea/�\�#Ƀ���RRݭ�d<�����X?WV̂BC�J3�.�� S}�����xx�y߅����xR�"|�{*v�E�6����N2��dM�$ "����:��u��p�'���1��Y���qI�n1�.��h��w]x�L�08aac��jh�ᔊa��߾��?���:5��@1;m�i������.���"Ǵ���v؟)wwwS3�UT�lX�"=P>/��������?,�0{�T�Pb���2Ƒ��O�\���ѱd����bQ����
)�������[���$�܉�sFRR^_�G9�L���P�U�����3׏����h}���pBt%-��;{{�1�p�בP͂�4�����H����& ��Ķ�@����丸ۀn�X�;`�4��b��7�XD$AUD�p�x�M�XՅ����9�<�a	"��A'��ǁ<r��}?5-MlӶ���X�����-��u�;�`��_����؁�gUh�P��3]6.�\��R��j5lF~���5��z,��W|�a� ��߿���F+�-;��8����^���l6�P�|�S���o���ȏ�)Ojv�0�Ǿ���R�?�w�(A����i�?�C�ʪ(��kB��<Q�����x���͛l����6���Hx�c��ꬼ���#��y�U:+��d�F���o����&��7�U��{�Y��Z���K@Z$3��l�f*Э�2캿%��a`�C��45�Q(����ƽi
"�q_ޕ�͊�ꀽ`��.������2O��m,�;�S�V���uB&�/�rr��Vb�� >~���]?M�� rwqa/ 0,l�wL�C������\��Ύ=�3B�{R�|zȱ�/��2y8���մ�	��ǏHV�¦��3 ����kH�ap�)����������M��#/�Ў�! #T�?;_+�?�lD�l�ϟ�Z��W�p��'� ���a]�K浹i�j�!zQ��
֛Ӑ&�_��ؿ�玦]��WLj`z�`��G�R�񉈒�x*R�Ӄ"�># �ɑ��	��M���g�n,�.Όc���wE����'e�)����W��d(��b�z�}��(���*\WG˅}��¥#��ޡ�DEC�c�o&d�f�p�<ic�-�H��GD�e�JK�
�Ջ��*�X��r��x�?%��A��q����X��4@A�_7�x����F5�>����j��zoo���M<��0�ѡ�4a���s�;� ��TE�s�~�%gF����嫕�9�W�)E�>m5a�� �Z�?�͞q��ox��w�޾��Tm�E�����2@4����򛛙�N?���Ȣ>���ߦxF49'���g�W���,��z|����܍�^���D�ʂ�A�}şLsFMC���������D�ɩ�?���OR7/a���n��w~JNSQ�ӛ������$3�XTto����ӌ "Y�Mi��a[�H�r�A���9?"����cz]�()���8�{��P�?#8�.]��|�-:���qI�a�W�����x �_%m!Ԋo���<�7>r���=�`1j���ʳg3ݨ+�| m�h����=�x�+�X�0=͑X�~m$�y�n�A�׸)V����ak?���HF���R�80�v�Z@�׻���v���J,Ǚ+�T"�	����E^��&� �x�Q[AA��桎��A[=��4@��W&�-�-�sssw���ц�o����\Y��(��9��ɓ��-lШ;]����I�z�Q�f�v+Øm w�mR�nx�2\�%%��͝��x���(�ϛ��5����v80�J!���c S���Zf�	N�z�o��ō Fi0��5m|i1w�0���dX��;���ɢ�}��S���D�1@�����Ǔ�?����,U���ٳ�!�;Ċo�Śv�2��EXh��"� ����;���zZ1_`#�;�Gϗ���}��x4 XZ��	x���50ͤB젍�?���-l�;�|Ά�z��Q��C���h}IK����8�q� @���FHXq�^��t$�oٺ�z�ϐ��I� �e�6q�<��<�jg�'O>.];/ݩ�XA�֪jw�{=��5�l�*�?C�,��C�p-@Q�5������~<���Viԋ�r�v��K4r1|�Xh�s{��CZf� �8"�_���@?T��˱
M�L�$���&֔�������rv� ��,`�9�Z(�®Uoq�����H���}�_5���pa+���gAE"L�LHL��7M�w��"kG\���g�b�v�,ZH��o6�5@}�Ν3������������A� A�͆Ã�/���K6Ӭ�QSSϣP���f�wx��[O�W�Qȑ ���S�����Eg�]��H��ڏv�WM���=KSRvu���_�3֟��Nت��$�:2�p�.�!��o��tc,�[����"6�p������E.��P�\<�k���s�nIś��P1I�
��}ĊƂ� P@��f�Z��.�&����*	 � �y�=��Sc= -����@��w�e�ͳ��4����&ѥ+W�AL�(_R�﯀aH�>��GeT���Ӣ���x'�qR����MN��f��C��Yn��ː���:9�����z��y' 0��zV�^7�:���%ߙ^)�Cj�w�9���c�v�sk��s��WU�C.R_<���7.?L��{u5�'�}{nD���g�rox)x��������P�7�5�djk�~��Iք���܁K~b�����I�ϛ��5πL�88>:6��@��DW� 8�&9��)z�DFOHx8=U�I~*GgqQ�����p��������~��תh���ϟ���d��m
00���)ukcP���#""޾��^#&!�WV���J���?>i�v!�}����njC:f�0�M����l�z_2��`�^��O7��a���+������E�Bq��Q��Es�\�~ah�Zbb�ij���r�S>�wgިE���TU��H�5/�L�p�>qr����^��f���3Ʒ0j�T����\ķ\@���п$��x����Pa3�k���.�;��^�}Q�@Q����%��˭=$$^yyl�UM8��[[q��8R!�Z'޾{w��=/�ѫ��'���kS�l⩩�=�.LHx��.vW@@K�@km��OM�f)�98��KW+�pv��3��H���ҏ�����U@�r�22.�Lw��� �e�狃z��O������llO%+b"���,�#JQ�mX�E�:��[�O;%�	ܥ2+D�F��4ܡ���|�3t1>܎G�P�L}w ����RTB"��&De�$3d�U��{&�J6e����&+d���#{޶�u����������~_�9��z��\�,mx{�zr��IA��!K�u�ۣ���I<ve�b%@o~��b8���0U_O��֠�`΀�`���ܚm�袺u���~�N�c���e�w��Jv��m�(=�7���;_�(G4g��h'�n�V�glԹ������=|5�;u�}7����ݰ�[��$�������L	��E�gT����d���77-#���坍��la�Gu��>{�qNAY9����ˏ�1E����ca��g^l	6L�Q�U�R�k�~�/}h���a_iPFj�&P:zܟ~W=�ބlO�l}專����tA����S�UTZ�хy떐���O��)�1����F��!11)�8��\ g�͛7�R�D��n�����k�����k �)?9|�Ǚ��n^
�`F&��X� �8i��Ű�	��ImH=N�k���d�Nn��, or�U�p���c5㝺�-K�TuL�dqQ�T�'�\�MW��Jr�~�I�Am5$������#�_/M������Wn��pS��>\�GL=��
_Sȷ_S3��`� ^�P_@!U�'�~�$�$H0�{(�K�.��9��/|���XY�Ӭ�Od(fr>��Z\S����E[[[���N`	�!9��ĵ����)2��.�1<U\�ǚD�i�0_�f��*�r-�ͷx^J�}�쟟��C��nWCn4��(+WPL���5)
�ݥ�3�$#!Q�=�ϞV��BϽ�N������Km�\�S(�<<l��oD�pTUU��ݹ����,Q��x [~XDlG
	�%J��'X��sx_���l��̸�����1M���mk�~f**a�e#����%=z�Ʀ�����bi�E�4���j�Yj��]J�M�,--5�:�y���J���e�������U�e.ґ�?-����F�)(��x�ot�Q��:��IEE
�{��b�3m.i��%eW<[=`�x9-ap�K�	Pkتh��(�-�VZ,f$28��0�u��p�[�pӰ6<�.J}i��}��;zRo�<�i�c����j�Fg���_��G	Ga�0$W E���5i\tᢘ��&�z�ϟt/sKG�,+�)&��xx^ھ:����Z���?Uf-���u�F�
 �b��~���C66E�X�������M}��3226��NP|��"5� U�n��2h�9��^m]92�;��  ���2s]��HN\�Wuc�63��䖌z��\��ess�xb<<o����]:�6��6�Q�*R�ih`Ç����a��!���릋4JJ�&.�J�S�u�X\�ɽ00H�5�Ǐ�}�i����y��ǹ�ۘ�m�=s��
����!ûuM�mOq��Q������[�d;_����D"S,ioAKY��F������R]��q�zò"<�b��OOGƔ��_�e!L�ˤfc��dT�u�k��~���
���mX�&#�lH��	u�f9�z�\�j8���|=��y�|秈K�"�?�O� #)!�څ2�.�!aQVrp�b.A�1̣�Ly�N�}���@?����s8	��߬�<��	t��-V�A �xx�����֙�K�iָr�y�6E/��^!b���hg{{ʒ�{���g"�|7������33#G��
R�3� BF�`�b':`7��K��s�\s�X��?�-dj�Է��j�9BD7��ld�?�6HGGG��dA�	7��+�r��OF 01�bww���J/)vtL�����b����`��/\���
篫���>d��vwC��.e��cʻf�5n�6�7ǂ��@�f��ճ�_����h�j2jʮ�� ֶ��7���+w�>7?/ޮd�1Q-�c��uee07>3r�/����t��%^+(P�md��m|�ae�0�K+lE������7���������/�.&�ԇP���2v����`�"w�������#�b�p�3L�NM鼊�T���ĭ�����d:�����O��4�I���/S]t�..)���UU��{���!\����U�WK�F�
�����b\�1������3ӄx�w,,����"Pbc:b#"�y�?�IH���f�n�'�����N��1�L��i^J�loP��Ź��S���~|vx.*@����RхOw��`���mz5f��J�8e����s6�1.Yn�H��u_JJ*�]���+�����dL��TX��#��ts]سe�^��_�>�''�,�7 �����Y�}}o�F����{�y}�UyNF�:aGHB"��M�j�SQQa���
k 23�78�1oߞ��nq�=�L����֤\�}țk�l�c��x�ztt�<���?I��ʈ+��u�D��Ru���D<%
�#*��)]�wv�f���$��>���Mo�����u���n���Y���?6���Y�R)G��ir�QO�e�
������<�n�
8�S:^�X����7�@���#�R��Y�ȹ���q�c6�BBE��������HIք���]5�>�ܵ�~�d��� �h��Ͽ5������+����ޥ�>=�{���`�f���B���ϟ?��f�o�m��o"*��'��f9�l�FGż�Xh�R+�;�mgHnEe����' z�.�o�܇�j�yLJ'��#ަD��aҭts,6���t�}�����>��[ ��331\��M�)��ż��5�����C�ax�x�\LI~/HK�:@(���1%�z��l%�o9\����ï�~:')#C���UQ�&�ǩ���gNN�L�N�Zw�	�& �_� Ac�^T���#�����U(&��G���>�j�m��i�$K$/��Y�W?�5u������Zļ��7o(����G=O��x)�u<ksQ�����c�3��xE
����/�e�(���jmm����|EV���XbN�mlRX˘5+�����o�����C&D8��F�m���t�~! ��Ȍט�:���zW�T$'�t|0/�h��$>�����/���N�Nwu�Օc�%~����R�x��]0�@����s��g|<�]���҆ �;_��y9XY�@������*�]J��oYXV6$�4�_�ʑ0����ML�fl�ss���g�������ฅ��!�;�ӄ�N���w����b�ff��o)���?��"�з��6���S��|��K(��?SK�������s�8�#E����T�Zf�f��I�.���H�!�>QlB ���5R��������%������#����ԲO��rNH`��{z(����X�����w ��o���捛+W}Ғ΢�%>w���p�OD��8�����7z��.���LT�;@8��v�V﫽���\L�!�Z��$~��Cv�,��U�/��ㇾ�f/;>�'��YR��n6��4��(��F`�Р�n�J6X�,�b	��Z�!��D�c^Jan�[g30�a�7����d�@a����~��U�>�'�

�3l�#S9�"ǂ���C�]kN�OӋ"���{�6��e�̯�q덮*���2��� +Tjݫ��w{8/�w��\��S���zu۽`����|���1Q��3��{���%$L����5^� ��Cκ:�M�-�hOמ��^��mJaY�W���md]�ʬ`�K�iT��<�bm���/����M=�S_��J����B=\�n��Di������3l�G:�	��_o�j�7=���u����9�����������* ��n�(-�9����Z@5&*ڋ��A@�>΁��F~�՘W�$쉮����܉��wC�2�s�cc��OcZD%3��hQ�����q��z��W�G����/p������>��t�A��hu'#WO��_RP�^2�-�l��}��o�*�� ��Ζ��߰��ܫe��������۝�JY%%*���O �Q�Ȑ��G���kw�O?��ןhȃG�a�,m^`������{����U�[�yo[��]WX�෾n������L�ϗu4WQ!�R��uH����V-4o�玣���f��23���ӌ�0�E�C`�j%����ɮ�7o��8�������=�8ix��FC�h�?�224�&D�צr�_Oϋ�gsw�*�����'x�p�֭P�pDsC�e���}�7�+0�jCg�%�Qo~n�{bbC�P����C��W�q��}Y���;0NE%j�ϝP )&}c�e o~k���g�("/������7n�³Q�u~:y�T�ߞ�ۈ��홏���-w�	�܋p�z���`#���fo��Ȩ�F�B������|������u�'o��u��x�O�H�u:�e'���7H��Z˕���K��(³�"�u�)��J�R���y�󪀐�2�J�N'J�G�,"��#<�j�r�����b�_%��Z<��(�ذ��j�*	{U���x�'-t�pZQ��˧�g�����I�����{�H旟��ޫ'Է�Q��X���=�bT���8wєzgq�-<)����^3��S��	�ttu�ȫ�)��z����潠%%&�ۿ��\��\���k��zJx��ϟ�Q�Z&V* ������k����'lR�I1�@|����*b�>�����y�ݿ���4����5��W^�^�+�%����e
�cA{w,X�1�W��6x����C�""��j�cx�?w��d�g�6C�C�WKF[9	��Z �[�����@&�P`�D�U��t���-G F����F6i�z�%�����a%�b�6�&
���Ӊ���-��GF�l��������11E��=��<��hSJ^��HF�
��N�r�0q��OTTT:=�/�
��9�wvR� �)(x
ܰ*�I�@x�-;%�::6ix���p��E'z���E���7���]-�,D�l�P;��E$�g^��ػ޾��㻙99����k��vu��l,T��,���ݧ�fӑ��v)8�QVޫ��ۑ-�P\s�P���/�|]��~)��J�F����/�.����4�rS�rxJ���aQ1�ay���H�	|T@����^6-b�T�D�1�}l���EʓGO���;m�cm�D�j����F��yX�(f����N���	u�UʌB|��å-�vh���ba��י��j����9��Y����K+@�IV}�|uU��@|���&W����j#x�I�����g�u�:)!y��H!��55r�c�A(xc"b�i�ro������V�?��x,�wԔ���k��O�Kk����:D�^U8I�p��⧏u2l���p�a��j�DDB�������}I�	ВF�Dw[�������f2x��:�j��&���N�4-�`�@	�>����+���N�)B���i�&��j!��0�ћ>������acb�49{��]W��ח�͉��OS��bg,���vT��IJI�����������>���'p��A��1T�S�SrU�;||J��8����՗p��\{��i�t8�
`��4�w�!�^o$N��j
+��_������7�"���nt=�sr��1~�:��,%%��ȗ�l�zO��h�qqq��y���& ��2w�ū�W�L�V@���a񤵮��p������K���z-���-�K���~��Z�������$@�)�Z(�dU���.��nFU#�J�|�#J����-�Z[;���9�j�{�6;�Y{�I@0:�t���'�DA���'���ƾU�ʷڭ�5��p"�����U��F���ǥ��c�!"zT�Hq�5p��k���'�k:�/޿�����I۝f���&��3����!\R� ^v�Vs������Up���'�
֦���--�[��X���.������W'���<N��V�G�4ǣ�)�j��"�
of��8��!
��#k�H�A3G��?Na4R�R1�Ϝd���p�.���o:f��$T�o��Ɂ3Qc1�O�yG�SX���3$��N5���@�}��㶻�LeBL�+�l��;%��@l^y��y�����o�{t����;K6S��҃)�߱oܴLM�����\\��>�� ߓ����ڪ�v����d���څ���kM^��F.�f���e�KJf`�:�I���5�Ç���$Й�x,[)3�����hs��$�ū����X��l �q|!�ޝ�g�<�Y�x���l?:�����J|�����<�g/�P(�t���໹{v���}�{�	,��':����a:F��h��K�)��:,��V.q;��/gP�	�P�(l�x���y0O��ܠ��]��j�9����Ҕ��:�F*(*N�՗+���j��[��I����~�|���s�٫^h%���ӏ��Tѻ��xI���&_ji�J�q�GYtW��Ƭ�]:P��<���~f�-L��JQV����x)x~��EY���^�ќ]:�w��S,'g7�ڧҪ�n���\�s�m���I�h��])GÏI�dJR�(4oĕ��RR��@"4nͶ|��a�E��	�փ�|�������LCC&'S��mh�s���N�����r�+�����q��]\�|�i���U|��Q��w\/�_;?����^o~@�)��%��r@d�Z�R���A�+�oX�#�X���H!C��YQ�f�A\�6/%���444tt��C !����>3���;�M��o[�����Lťk*�b 1Qh�Q"��;::��MS3.o!������+�-���[`Q� ��-���s9�z� 1�����R̗s��$�c`���]1�m����9=F��"��{��������}D_w��J�55�DC�_�F�jO�-��cAs��۷R�1q Xo�ӊ�3w�oO644��:)�)�����P3�������#Œß8Q��龗�==������	a�Y�����l��=��Dmx�v��d
] �Z��B����ş+�Wr*�
U��{'�2Y��' �����K���&22��g]UN;�����(0�8�:s��3�����́sa2ދW�s����{י���l��ū��&Cu+�
��"�ACG�UV�� e1�%))	,�榥��������o �����`S��R��<��� b�13#CB%��? �#[�v���N��kx��e=zz��ǹ����d-Y˗/���{r2���~�K�!+յ��-1 +ˬfY��*$����:�9� �8��55��9
>#
JQQ��9Ccc!�{��l�jjj0��n���n�A}���1��MllQ�������mo��;Y<��jF8=p
������+ \�	Ÿ�6��B�oe�m�G^��9��>��uW42�B���@��|�Ȏ���q量�&�F��-�� X#v0�o=n.�%$�a��0Ĭ+_і��2/�����t�kc}]�ͭzs�+�ˆ��{�� 2�����376~qF�x9�����H|(�!a�� ��db8A4FkiBTTڑ��G�͢��r�?�*"6�3�����F!�� h��F@l�E5��X����v^}���%�%p^��_�	����� ���˃LC��y��K��z��	�eV������f�����g�z��Byt,lؔ�W�O�^�]z\��q �^��{9�,�g�6x��ʢ�A��|�=�����zsQ�+.*���q���l��b�7j�-��@��Iy��d�`I0�Ϥ�=�E���\Xl=}���,Ѓ��)(w��x����T����(,���*7�E"筗�<O-�lfj�J���{���'�h�-�dK����6�|���m?41��9��Z�&�����'rq����Q��ˣ�{�OJG�J��,z?��M~�݉)�L�x}�g]&&&}�FB h!�}��t��������'�Z�� ��@�7��uq�����! �4�-����W��Y��I����ii1z��N��I��5l��@lhi���M^��u�JYEEj���E��=%����+**6A�n}�%�,�]�`<�~lF���Sa'N���	��խ:�������~ \ʒ�����b�kj�a��"�	,cz���H�����/"$0��t� s���CmcL�=�n���Ds��!	l:�tl��A�u�x��p�isT�.�t�r��G�RVa��	��O���e�33��{G{��]�/�҈?��F�o``��}��,�636�/�7������CC���lL��
Z}����]𫫫)$���d��Ʃ��6�	�8>�J����c�1����I�k^��u//��J�c~^�߿ƺ�x&�2��̀�����h�Z"_����ʉ*k9���y(l�������Aڣ�x�x�no�x�d�+}}j�x^��O�z4��H�vvl�;R���g{�N���MO�{5�<%
T)6�ǈ\UV�i�&S��xu8��D������amTE�|<<�*��~G.s� [.u��jseJ�Z�f�%7�.o�guٔk\P�ţҚ�m<���x��X��$�,�vw߁'��	�4�8���*�O�(A>�f��w��ϷuU�z��@ZX0�u�	3��]yY�c��O��J���W��z v�����~��(ld������ p��ٸ�V��Ǔ珋?�˧:�i�4CEEu\/_�엗�/���U"�u�qe0��E:���-qaQ���;0�3P��p�Ľ�=���r�p��ߝ�����h��+C�Q���.�{l��b��II�r���Y�}2�Ta���XWxd$�e��Q4�C�<���H0X�O�j_�@�	Nhʧ-
�(�������)S�[��	��$e�Y�m��>���㴺
Tf\5 ���5B��-�j?ss��A [�K�7^�؀ڤ$��V�p���c�u8�]���xi�����.�/� 2�3#��ކ�m��[	Ę�!Ll���X�6�&��@�,��5�2����#4�o��ҳ���:M�Ƙ;����e^��.h�P����:�QQ%^(�Mǜ�6L]]]@��}k���_��k�����8��%��p�"�FB�Zż��}������d�\ �>1�����Tg�[MS��-�6�H#�������_�_b)q�u}�е��Ɛ��l��,�^ݸ�k��c(�0�~��#`��ջ����M��8<c�/-*�3�,&�:��V�O��O7ס�P �B�?&i]����Ba����F��.P�F[3MYP[�A&W�6lU��$�^�̐ŵ�ɚ�V��->gk/���V�^�����ⶶ���?������[�ÒÝ�X,�x�}��~v�1����@�\������tZV6aש.l��K�io�v�>�e#����	P.Rϔ�ը͞����)���n-�D7�����^6�f?�p+��N��[�`�5�1q�|r���N���Al�V���aE�4�K���,m� �v ������������ݗG���� �x��m�"M/�-t�z���'4�奤d����H@o˷~h �h�n�$�sV0~P__�Rb��"��,%�{{i�qŅ��)e��@��Ra�n���7���R�b�_��d�6��u���b�6����l�hx�����"1�_���z��)ҟ]��� �n��yj�@�$''����y�}���3^YZ��f�w�oĽ���� 6(,�o����~�	�{R��}�`�k��RŸ��D��3i��Ħ~"�+R��1c����ޝ1IYY��鿲�����1Q��{�"T���f���|�Tđ���*,�ޚu]���>P<l�������Kp���u�ن"����9X
����Eaa<�piˍ�5���k�q�M��* ���1111A9�^���R�uk,�ek�.�P�˅u�r_�M�c�N�t\RZ�hcF�2�i��1pU��~�k�ݚ��c�3�jU1WS�2�qJ�Υ�zx'dCMMms�m� ��ݳ���e���.N殢��b�*<�k�!�q�!���_�	�\�Z�0;�}����L�����T��F�؟jK���`��z�R~>:2::q��@Dg��-`�T+�����랼�>�ʦ��Oxi�amCC���S��e����c]���),�k.��*g�/P������)D�<z�V�jno464���N'�"�6<Ώ��X�8����i#����"����///׃�O�IH�5�L���Y��=w���x�<�j緜z_d�7u|�nӼ���N���e�StYZZ��D���[l�{JN'6�cq��)&_�[f���q,�5���и�����\#EEE�?_C=`�(4$<��}?A~}�7�y/Pummmgn��yy����*�(ie��}�i�xzU�Ɩ����W4����`�Rx��躑���ܚ�G�An�|�/w,�Za��~2Kv���S��yxD�t~),P�G��7Gz%U5�����i2s󜙷ɢ^�H�;�� ���Q6~��imf&&�l�b�aU��
PS�oR�C���KG���s*E��|\���}�$#�[DDJYH�2�����-�M��>�$e���J�_\܉N����:h�#I�C=W���+�zmK��L|x���%3�����o���o�̚��ܘ�U{h����w(��Ȩ^�}�UXЍ�Z��oz�M%�W���X
���`A �8��� ���{��P�L��jCVv�ߏ�|s ����[�n�NNN�d"h� ,N��O�I]7��ݻ��x���$p�IH������$�'E
�;��cPP���럱�t*��o����6���\@3}L�:Ě���b�U5l���t���&��"�sA%�}q�v����r�cL'?���?��34$���ݸ�V{���U~w��i��A��eG -��Jղg�h7W�Ϗ2�OD����M�+�!'=Ύkω���2��a
"��<������(�=##0]��w�ebf�oh���LJV^�Y�sn,������vl�I����4�����5::�2��o�6S��cFc6f*e���� ��셮a�Ê��q�^w<���<�+�M�#�v�B�f%��vR�6�;LF��8p��ۊ�9��:�S�Zj��w4�}W����v�:�u� ����dg�0���%�1�NŘ[Q���"S�qhS/4�<;�=r�)���J����l���V|�Ǐ����211��$+�CDD$r�M��YZ[�ɐ�� �D�@����ZR��tY��~����ëҀ�>���461��e���?�0KXW�����/����=�5�S�yx�
{�]U՘�Ö�������H)V5<���1g�q�yL���Za���Du4��W�<�Q�
�<�h21�{>�̬J|�q(EK��v�nw�/$2�0�&����6n;O_�*X�۶�8y�e���t�_������Th��c�]3Ě=d*�J�wHHJZ5br�h��o(�o���l�Q��+	�d��LM�$��TL�e.]����f���XVq���%�N��El��R�㜧�f[��(��===�����,~���~�/�-M��4UhԔH�d�+�gJOO����0�'��&�m$�����1����ȥ����tFᤈ�5@��f������CBC?���ږsp��}f�À���\Gɳ�i�\�G�ڹX➓E˗���&#��>�塥���0QSV&������TvΠ�o�����������"nǼ��o�v���f�w��j �����(�y����i+�b�u����aw�Ȃ~����BI5��������y��w�m�"XȞ��,���/|6������RD�<<jg�������߿������3«��[aI�����mmYuX�p�߿���8M�����=4�����k�VWW/���tw�/t܇�ȩ�o��Y�����j�D@S F��&������)�^d������h���\�ɲ��������x�ˤ�F�1q���7�P!���/_��Р�˟��.+p@���\l�n��q5t%���X}����R�'�]	�p�z4
.F|����ܛA����'@`��>���-dq ����ӗffLD���(X9.k��\7����h󻵡��D�ll�m��Cո	�%�D' ^e�?;�����8��]X�CVV��c{�r�z������-�%7�� 0�͸<�����#e�}��F�!@��������F����Pݬ|�L���=96:����'�D$$r+�B��wQ
N�m�G̬�.����$�`�]�Wsv |�ϐ�'"7=���(��K�OضO�#��8�UL�:VÂ�nhh8,�wG`E��[���)mh�p_�]�&)11����ܣݣ�<��zϮT�VX3�qV�ౕY���}�D���LV?��o����^�?d5'�ϡ��V�d�/��F�U��D敫f=,�x�Db���<��E��d�����8ԉ�eK�֓��ʘ�N�m�	X�e1��-v�9��<�s�:?�|�t�Y�pO�3�\ ���lC��p{�q�ۻ�zt�Օ�b5&8Ь��/���v'#��j��L�ѩ�(,T�e�n*Wם̽}�����(���Y��^j�4�}1?�q ]��us��A���uy�sf�,�E)Ϧ⑍&:��c��.¿�jO���ǀO���so�07��,J \�&k��6���6ȓ��
�Y�i�Y�&��X;��jg��'������(����i	��ӓEiT»/��oKZ��9�M�f�|�*v<T�М�&����޷�muV�>n�z���EK�MOlƕaQ2��)#|���^V�@��6�㚍���p�_��*``D��b��oEm+���I��5��v��p��ҋv�}ظ?���ӆ�n��om��y��v&��f%�Z]]��R'�\��	P�⹘ugm��4�����+�Sz�I8�F�N�mX:�=
8�<� ����$l����6obv����[p��%��]�{�k�p1�Y�%2���qC�Е�,^��׼W�R�#���ݻ�:�R�^����;����Z�R=n*�j�X���D��	�����U8bi�5�]=�;�~~��W8c+Y��#M�5�۬e� =��ބS�9��Ӯ䩘f��`-lN�EFJ����P$B gW����V7��Sa��!`�15�E՞��դ�{�$R��\�w�5��tnN�hmD5�imT�>��t))(gi%@a0��.:!�y>���3\X�CpzT�e4Zb� �֢�O<T��X�K��Dʌ��#X���h�.�
�r���o�L��L��k�#x6��O�2��]o41.�\��&�HCv�`6H��z\�ƾ��a�[\:f-9�0����Ó9��o��l��妥���>׽��k���R��+*p$�FQ`����R�aޘ����ϨwS�(����hPw�S����b�����$Q`�|�1؞}1Q+S�ő�_mF�n&�j�;�J�I�n
��b5�U�u|����N�q}带vW��'�S[dE����r��b6�P�s36�x/�c1�:[����N�&Sq��|
]`ik���!��F��7�� zԼ�	����cocc�5f�Q��;�
���]�bq�M\����L���c4� 4\r�%<�ތV�����ua��ݻYĻ&�q��hH]�_������`-k,�6������=��Nl���x�2��ԓ��bRKL}F�o��οZ�Y�%c��tY��Y��c��#�6*Vr��G���7j`�R~)�l��Q���X�����Z�8�ujv%^���UZ������*�!��4�=�S�d7S/'�5��.˥�l6��ck��=;�u�t����5=\߼I,���OaJ��a�(؀��rv �g$M|"'+r˪ېu��6�p&?t`I��9hb޷J��Sſ�����0U��N�������ѐ���oI��a|����5���?��ø��ۂ� ���Wk��')T-�m,ϲZ����*�#/�w�m��}�PY�8a�'uѢ�W���崄��Vp	��	�58��h��@���t���	��gϞ��Xa�M.=b1�#�_�����'ª� ����[9�.�p�XN"��]f��;�����qs�I��'mK�ȴ�l~t8�%u����9���c��k_��{bv�������v6(�IzG��{���^.I=t`���K)�v�)�.��?�
y�Y����Ό�8�8?����>+���ϲd�v>R}��xc�z�jaW$���*'z���S�t����Q�l�����E\�i}�^�r��X��01�@��!8nᄺ��?����2���ǒ���;3K���_V����S�'�Z�=[��:C���������7�S��|�ˢ��f׉1F�߸86h��lܼ�,��7&������p.R��1�a�L�J��H���ROR�*�y<P��1����!�!��Q4��d������WW���J�+���L0��}9��]â����v:��j'%��X�|�}>-��촇��Q��d�Y�����kठ.ׅg����k� OY����"{=Y���/l�VQ��8[b>^/'j�o<�2a"�I]A�sS��%E����9+�u�>2�����ץ�&=��;��Y_M�o8�Ix�v�i;�Ě���f8��l���l)茎Y��t<������K��2I�ڠ2ȴF���^F�����?P�����i�Qv��r�/tK ���[MO��Īب/Un�mG
jJ_,�O��(�{�w�Y?(�����<��d��v��1���ʽK1h�#=u|�<r�.MWx��������s��̇������{GlA�2�TH��S�t�ߤWr����`�t�܄��䄋m���~m�2kh�	�·���*,��`}Xb"�_?K�8#�X{�7���pCN�)AדY��]c62p�x��"��+�T� ��kN�V-�AY��� B�t�2��ɿ�e3��z�K}f���(�h6�7 *�]�\�vť�Z.��w��]L+�F����ۯ��/׃#�*k�+�GŢ������Z;E��G�%�\�
;c8�|S�8p:�/8��?� YM����Mn�P@�R���>a���MV���u|R+/O���7&+M"���w	�Ty~��,{�հ3:�-
*�_^^�>�Ώ�(��eɾ����x>bH&���-����`.���A�����E�9&�|r�:�d:��Ur`9��XC���j&�ɌH�F|K����/��6�܋�Mޯ�b���E �ʤ^�+���`��������H���I���6��徴�l��\�>4��qs�����i���^���6��Yd�삣�. �����|�f�i �s������\k�ǥ�G{+sp�+c�Үh .�����1���c��"~^������Ͳ>�����+�/F��Cv-�AO��y����3�ܦ�^���B�L�E��n�?y�6�E"En���bz�Ռ0���@8t ��Y�'D���B�g�x���'��j�,�����ؾ�U���œ�2�t3����	�я�b��*����͹c+ٳ���~(�ߍ�U`nI����T�3�wZ�<xT\�\֊�����N��ë*Y�i��7$#K��ͱ5m�
vUhe���>�y�����ut����%#W��?��n�Ц�	߾�Bu�1��3oKg��HA��trR��:�$���Ы��'H���D��� �!�s�i�y�*�ǿ (�&E%�ǩhT9�>Q���H����.�}B���J1ZR��r� r�|��m�ժ&��R�9첡��4�	U2�=SXCН{)�u�{3��3t]�E(��XТb�$��w>����	~��>�f�H����dw��^��Y�C*�OPXl!�(h!$L:�+���ܑ��O�9�o�4 8&����I����{��Փ�v�.����<���s�^�/D�ْQs��{=��[-d�.�'��R��r����� O�m	��C�\���o��>:U������4�����O��8"�[�m����sw8$|��
�$�J�/�%k�-�[,�z1��7�u:��������W�����F�����a!�oR����{��S�?	dpT����3cDR�/��p��uum�7�h0���3��M��H��Q�ON�'�G
�ܐ���0�@��\c�Cb��>`�o-�#�(�ﲓ�Jr����"�J|׹lPI���w�V.��9����'�����.��ow9�})�4�mZ�����]�K��5��!g��-`+_KG�+�/,,�@B�����d���U^�[����&Y��Z =��kn��5>�υ!liE"�0E����z�D�X-lo��]>}whu�f��<{�'����DV)x[B?H� $��Z����I=BR���ɚpIU#1O�4�A(�׽T<�@�p\%�l�����ɽ��/|��|����A��H]V��BO�5�f�꽬 G-h�" ���V:��i��<��M�BXl3�0����:�� A9�1����}��|(�EC4�3�����`x�>���'1�^���j���F�-=���u@޿Q�t��?X ����ws[�d���>9L�\��|�C��fG��2n}�&����j*����\#�K�ŧm/8 <o�F4��4Wӑ��U�[��C��X�dÎ��{�� �w��޳׸���F���(%` ��&��߀.�q�������U��8�z4g/mv�z�dk�l�6��mE=�ac�����RJ����%��Ó!��^g9W��%W�vc�z���O�|����b0����(/��l�r� '�}�ڬp�hg1��n�T+�5�����0J)�c�K��~%2l1Cv��w��q��5&���J磾*>�Ը|�^dɸ����S6�ƀ�1OڴA��+D�����!�y2Ej5�KJ46}H�^J�M��j�j@|&�Y���e�����dv㴺���(̓�b�G������x����o��p>���:O�K�S)�N� ��5L�N�����a��I���;��{!uB��G봁D_�� @��eP����]ӢJ��Kp�\��}'p�z9��у�|����b<js��n�p�Ť/�/X��8�H����a`�u��mP��d����X���?6E�e�q�Xd���� �ƣ���zͺ,��(��$"�e�%TS?LHV%q^�s��A.�޾X�)�N�m��l�L8u�Y�8>1���@b�f���	8��m�'�|8�������&�8�@�
�_��?NP�6Z�2y����K�����.��v�l'E�ѱ�[�\\�k�:�;k�N�>[�w��sz�UkJ�V�0�qph�i�f��e�d_��M�^�@��?M�6�o�V�8�X^^�����*�R���kΦmq�1��Vq�\�끵���r �'X�����d0фHb�
@E�fО����P���/a����@X�H�1����^����qs�u���:ϋ����3,U��ޞ��C�
ʌ���Kԉ�F�.���8�̂�5��ܻ�9����$ ��:���P�������՞�`;_3��4����l�8�t���Kz���oA��[0U��UL���;�{ O�z� ��ۏ��5UL$�b����G�k�����:	u�]��=����f�3��ϫ�-���U�v�t�����G��#LEB�4"s^�(��]�0�yn-/�*( [�>G=�H����߳P�C� Mh'}�t��y�G�x�fX��?
L^�8��YZQ��O�Odbd�k����3�Gs�V?�2��{=��c���O�b����s��K�1����nCV
�m�%4���ǜe2�ߺ�λ���'PK����\�Y����]_��.G�n��f+�B��ޥr�п�o߼I�n�S��rcgi*��\ͬ��������{�P*?�j-��r��������(�u�b��;\�	4$#>�e���ɛ6���k���|k#�z
u�򕼌�r�V��	Sv�\�),���CS�"�����چ�vn���E(C�&>tt�Z�'r%,<�Y�y���L��gS5�g�_Y_e��?(Z�Y[Ȓ,!��Œ�d�.��{fl�E!2B�$�"c�B�A�mF֑���޾���u�uU<�9�����~Ι'5�|^�����X�$_|�;yK|����t*7��c2a�z���@xY/̱�Nn�ߋ�hܼ�F�0,,�����1I{��`�b��l��	lC������JſcMUQ|��AF�g�ɟG��Aё����oAR�9���n�a�ֺ���\"	�W����& ����h,����(��p�p�⴨~Ďꣿc����H)bS��-1�]x�;� j�J����S�ɝ�]l䙢Zi�Ϻ�w§M�}�bit���b�5��d��~�x�z��<b�a}!M��� �!���ٕ�;���W������+�_|6Bp>S���	,�3#�.���D]7���м�����U�d��`�,��%�����TL��Jg�hFJ�d���E��dw}!���ls�0�j�<�Mlz}�����8�&�����	�崶�:�D䞞��?i�m����'n�y2�{�e��j�����{�=Ī���W�"�M�l��7Z�����ܟ���*����L��I'�Nt�+����R�N������];;�#i��4P�4���Z/�*V�=O����E����n�49R�k0�1�D���o����R���"��C'*�;xt�GU01�2O��Ŕ�~�����K9^^^]$_�z���N�o
1����{
ً8pn���X�"1���~��X�w=�7���`��Zb&�ӻаX������t�'������Q�y���|#Qy�{f���[��ÿ�`�VIx��`n��,M��5�j�4�`�t���{yU�U�z��]C=�� eK�����u9�~�� 	{b��5Yڵa{m�)�F("��p��d_����d$��+��י��J�����W$�$#�h�>D	�:[�^y3�o8J��y�3����Pc蛔x-�LGh��];�!Oә���zJs:�
w�dӯ*y=B � `Y��L��o�q>y=O��vN�\D�� ��YX@��L�'��t��.%O�����t� ����"ybm$��f���N�w�=!���h�����빳�yy_�� C�$����H�)�(�2��F����uyy �6�=���=Z8�5��@��&�B�,~1�5�nskQ�
�_�7��R�6�#i��Q%�a�u�o27�-��{ibڷ�&V�Z�Ѐ�6I��U ���N����p�^�ʸ��:��B*��\�2�:d�)�������ۦ�#�����,��oX5i8	�1��+�~��F���?J��%����J�H{����Yθn�z��$ɤӲ,���@����_�Ov9�[��^�K���fN\=ow%�9Eډuu�BA�r��C_�Wj�9inw��;����P���F)���m�@ձ�S R��a����5���Y���9�-�c:;�:�잻�۽�a�c	���y?�׺�WP.
���:)u�Y
Ҕ�F8�Qq��X��/xTw��l�k�󨩿ާb@�J�������1�A�w��P�r��{�(ŭO���;���g���p��!E���pF�'/E ���7	���F�kGƘ=1�lo"V�Tמ?Pu����P2 L�R"��v��a�b|
zQ1��O��<��� WXN��@��t
z��\w��c�k���W[>�ugA�uI��,�����w,̰�)/�!���BD_>_��_�W���vk�����x��-B��f��;�ݝ��F A��<��0�Lj�L{��A2���{�����5���͕������/7���ef&/��}�p�����޲�h����#����W�?q�7���X�7�˳q��p/��4�X��6U8��@�晻�i�G^�^��>o�h�&(��X\O�;@G��?%L#%�����=�X�d���UE��mѦ���š���L�C�����ؿN�(@x������:�+e�(I���<v�)-��m<f����s�C< ~D����=1|1)W�Q<sFE`�#]�qY8�t�~�}[a���ֶ���:Z�O�lw."MA��SSE����ERZ�j�[(�W���3�w��������:6Y�LX �@���B �Ca+m�����W�RZ�*��YXn�;z������镡���Z�[a�������U������7T�t�U����V<-ť%G#����K���	'�����a����NCw��R�֠�P�n |�ꟺD���x�l	��3/B�?���[�p��F�2��W�~�����|u|rD)c"��� Qj�n%�<���֧�Z��gs�� z9��%�O��
X��K͈N�=aK�/���l�l����7d�9a���$��PL����������x�m���������
�aj�5�d WD�+5ˇ���>vC���&��HJ���I���x�s'q��?��-���&c~b�RS{=��>�ԑ�G�yk�J�=E�)��w�&?��.:4}}�𚚐?�p�7p�^��i��"��(|��wv.��'�;y�ޣ�����ȴ�R;�F���UA�i������4I�L�or�(}��E���%��e1���d.Ö�����T�����tb�5�>��卮*�
����i��q�]j������^��p����s��GzZABb�+����H�z�_���IkOt�i�\Z�]0+�LP���'?���y����ެ����1�|;ZV�t���cI��������^1��3�㪝ң�%%�	�{Q4[��c(D)��)�!�^��*�S��7��w�x��׶�:���<�� �o����bw�c5��@�~�������Q��2���M��R��xO�IE�`K�X	��_�?A�ܔ�����*���ǘ���(�_��g��9�P�a�.9E�I��o:���W� �'���i-]).��Q���2���/��nwk�X9�]����_�ނ>��pE����}_�d��b�:���9#���`��$c�����<��l����n���Ũ��[#aU�7/*�T�sV?���b^e�6@�q6Xf�Hg/����ޗ����z:���!�A5sz6tp�����]�5��?������m%�Ш+W~odr��B��U�F��Ș�I�1�����wo�^��z�zBFlc�h!r⛋,�� �,1���\_�e�
�����j�H�5����Va�j���ޘ�M�]W�Y��PCxx���~Ê�̑����w�{�������t��$������|�9�
�-�RV_]�0�o���
��RbM�:Mu�}G����%�>��o�0?RkRsv;FF�FGS��g����5���ya����3��\�3�Y��������x���=\\u�@U�S�?��1<r�\��{�A&�D�ZD��N.��ԀM,,:�cz�����A?���0���7��[7j�{-kloA�\ϓoP��NQ(��-�.��n��v�4�<�����ʪ�ɴ>�
�	j^Z-�]�%���\��r�����+ұbE칽;����A�@ll�CG`�s��e�y�1����I��8`$����53��C�?�����X�j�ʄ�7!C���P�U�-f~ē�;��'Ϡ�6��
�x�q�TG�ĝ[\�����0��9D���ON+���hz�S����V���/�`7��?�1}����[��L��,�91J�g�����S{㰁�V��eիs��� �ir6����y�� �O��E�H�y�C�dΡ�U{t�<���&=,��9�s��Գ�hb;������H���o2���Ig&X���L�R���˗/�|���If�D~�����=!{�2��*a��\5ߞ4 f��)����B,
T$1[Mt]A(`�w�q,� ���d�m��0xP��j��M��+�a����N7�_ˌeț��셝N2Oi�!��dy��JƳ��g��7&Ѕ܉�u(#���l���z�hj��z�"G�8�3�g�v3��C�����p/�*n���X�h���c�n/��� `���c�L0�D����=3�w���X)�����?��7�-T0�-v	���r���[�:�M�Q7a�+e�j[���F�o�}����\ �U�xjYf)ův0���А�h8O��w��o�&�d`N5�D�}�*6E2�����(;i�ج��9��c�|5����+`�d������l��e�H���߲� R�h|���(��U���G{���3<h}�'����U�*`c���:(>����eF��=F���om������[�zT�K�`��0��a�N���k�$�J)� P�LQ�}���V�AŁݰu�6� ���]�D���7n��͟L�c�� ���0�g(�@�=-���YG���A�����Ⱦ�(���!�6���\6;���k3A�+�\WŐ�~U�kea	�t���+{����������(���YG5o�%f���xy2e���F���Q�\'a�Ϟպ�Sq���=" D����>���iy�.FVqA[Rp��:�˺��Tb�8��F.�d�G?:@�-��:e5E��i�?�K>��u��Zz$r�#/D�I1�ԋ���>y���?�������[I�1�[�����:��ұX��D�~��hd�uI!�����B�-�&D~L�ޭדCJ�M����iZT��P��/Jఙm�'�9�w3�����8��K5V"��Nσ���J�]������k�:E>wy=C�P����d;�V����܊��'{������%K��.��3��C�A��Zm�c1�3�ޮuK=�����^�.xw(�����АpW��i�$��1,N0-eC�P= ��V?��]�Zğ�V��\����8x�Y9:v������ 	��BAh���.��D�@�ϵ�w+��7R�v>��NP�{����[��U���t&��_E� ��Qg� ���Fa��������yR������!]��4�3�&$�2�:O���%�0���`�:Q�6���h](V��QA.sE#|c	^�����H��w&gq�P,��ܯ	�FB�k<ƃ3�g�� �؁X)H�e��E���>�L�2�4V��5
mY����c?{SC���[�y�	�]<���{�މ�Q2�`���'�xlx����B<��ܒ�����y� �&�xNx#䵔��V���`��\�T	R��9Rv�>�o�J����%:p���mn�W���]+��ߡ��c�����.������߁�9�,bTh^y��>\�6���d�4~�4un�)�d06�:���_V�x|b�i�tl�o���p�r�nS�f}_�݂�<bG�tK���)�<�>QEc!�����@_��;�C���<)WO�d�T���w�H�u��u{��0
Th��ZO��1LE�WT>=9Z�߁:ȁ�K�J��	LA�������!�;j����)':���	�F��	�
����呌}'<�W�D�`0u�c5:UYG!�l���p?���}K�Ch˔]�~h�e'�k�C�
b\��{`!q��qSo����)8�0���<b�30.,����%���6-U0�lA�{�> `:����� ���{��B ��g�0�梚{Ԋ��Cd��G��k��n.��W��l�c�:Ԧ����Sz��S'1�!F
��AI��T�$���b3s�X��1��@G�?������{հg�HD����}1���fsŻ�'�����T��� �Q��/l��wOXC&Y�u=E�w��iq��6]���:u��ϫ����Ȁz~�%���M��>-uV?5_/���N�M���2��.���x�k�������0؄;w�z+�{�˗O���4q�KF�yޑ��D���ص+k+|��HV1��t�f����z����0grF���qv����|��� /b�c�z�sz�`������r䱧 kK�u�?'���$w�=�:��}�n�E�y���%��4�'�-l���2�����o�0�v��݅����8�f
�
fV�9�lZ�U�
��:�P�< D�d-�z��|C�|@�j�G�٬�2�L�'��^�5��Ӯǋ�j{"�s�r!ch��2m֎k/���6��"�	^��ݚw��O����A����ð�_�_�}�j�u*��-P�?�{K�B7�}����������t�6:E�_.?��C�B�-�� qB�Z9��k��'77����0_�a�,FJ�H��?��M3jN2 q����&��
,�����j���V��k ��njw�����&�)���;t�K�Y��v��c9�+�BK�7W|��w��M���4U�_�I浾��"���i@(Mh[ϱ�;9�B�=�Y�m�P�Ձ���M�|�K?=S�)��.�8�ȷ��>�F�]F�6��/a��/����ӓ?��ʋ�̐�ʑH�ZlA�a3����A[��YZ�؞��ǦBug$��!-:�{��h���R�D=Hq��P�n�P�~�D���c^�����h1��f���r2."��������,�!*C���*4�=����BI��Y��&�W���9-����	����[�ƿ�b����rE��B'Ła/��1O�rT���5�_h�o)�VS}H��<�����9��E�u�9�$�L�S�-2�C<iQB�Fĝ���PH��������=4JL��()ijk'��q�]�.���tT�n��+��� �eP���9.��=�PT�n9��x�%$����7 �Ջ��j��[�죣��A�b�t�G:�os���"�!϶�1�:���"�?�a�o+�e�����:�9����#.�3|̝׼ݶ�3B�J�h��)�B���@��q�O�� _�/�~͵��k�~�%,PL���}m|r�� �T�c�@wL[���oL�4y��~�ε>R��Y�/��&��V�Z#�{	�Ы`��۝@5��&{RkP�Q�y�u�Ef�s뵊G�	��ͮ5UW����n� �n	��er$p��j)M;w�h1s-���6-���TR�Ѓ!-�d��[�4~�?u�~>��x"�S���������=�� �;�̗G�̠U������= N��˝�����y	(@�?�*M1X�������'w�r�LK��p�ӳ�l��r<�P|�>}�?9#�#�a��0�2��\�;-q�Z�#�C��p��CO�&-�@Q�K��Q��$ H����J@�5]�#�����O�-�m�[��S�T�{���P�uI��K�n:�S�Ǐj}�,�j c�æW�1�,_��3O��V�N����`A,��P_�;
����bC��Jy=���S�����%��2P<;�=�.�s��N����!`}�m�)��ݠ?���#��'������]�j豗����8֤�zS���Xn�=5���O�xq�z�4�<Ԧ�j8`�:�$��9V;M6��dy=�S�)����c�J
�fV,�s�,}/+��X/�S�[d-�s�,���s~G�B�:��
��(�<��e:m5�n5�c6g8���1k
��o�.oh`�O�Ί.DI;����Qcm��ש~�z�����1��zJ�oΆ}���S�֗�C�L��5��Pz`�������
:���������:����T����0���6Cυ:�ΌA'�����ד)���Ǐ��Q����'7��>Gȸ
Z�~���FdAUD�KB@�̕�F��U��>,mxB�A��)�c���x����U��Zw�!U(�U6)����CҞ,y�i��Y=8�R?�J�;��Xx��KV�7=��QX���g��s�C�� ���N�KJJB$��*0�9b&gp�I��NS�:�p~��f��-HRa�瑩!�Ѡ�֔9'}���Sz��ɿG.��g�_���������v�7Ξ�ZpFu}?@`�3��N���f�ù.����t��Sÿ;v���-_<�)ܻ_�?��ġ������7Zt��|�ʞ�������<�*�?�w(�>��2I�7�Փ���0���N��XD�������1O����[FG*u"ǹc�j*%k$K�4�YxZ&�����!�aCȧV�%����Ә�΀`�R�pP+o�r��؀�s���L���X�6������<r����ҫ��վ�b�b�)F���0�kl��]��:M�e�6x$���d�ӑ��x!5w�7��ۂ�H�z�u��b��f���F�z2�i���{�pJZ��37��@�U��ߐ��6���$�9��������a�cyO�ـ�-nF��}�Pl+��W��q�PrO����yF�&�	����%��
�0V�c�#��M�xn/ �7+&�W�4�c9X|N5����J��#ܩ�NXNٺ�;�=%Ȣ�鎛����;���z���F�,����tc���9ڬ̼� ��'�*����1龜��.���鲇WX;�R�v���}�2����k�u��}D��~'���}T5�KH��d���sd �?��y8ʼ�vk�D�6��i'}��_�2?xo.�P���A	���2�9Z�u�2��|�5%��b��g]��Z}��v��� A��K���[�LNm�c�jǓӴ1�P�`���,GW����`�K�e�`]Z�>ՙY�=�F�u�)�
$�'���_I�����\�[��s�%|�s�@�&���%�j�(�D�����*|7?��qF5����dL�]�>��@t�ǍYl���L~=��[D�;ۣj�{ʗo�;݋��P�EsC��������b2���sA��4�H���Y���X�x]` �B��X���$�$����w��"^��l���:��>bS� ����<���K�"� ���6��LkN.��������*�ث��a2wM��M�	Z���(#���|�w��e���ܣ���}8Λ��
N�l5�<���f�F��c(��O�Si��fP�O�h< {��̞3�C����pyyٓ�h(�-ȱ��E�E�z�\
��j��,E�*�r4�J���`��_opo�h���#.�W��?������Z)��*�R')���&�k�����`�׉5٘��خh�뚅z�����q6��:�9���W��#7X%X����j��xs�V��ሹ՚����u��YVÑ�B�#��3C��ؽ������\'|�f��0��L�m	��	�=R�� ��1���Ǭ�r
���5��S�z]ѽ���r(�Ml��"+ە�����"vM��	h���p���8���N��҅�;/_�����Bp���N�֧k�B0h��:������*k{�����z�BrOzD��}Mcr_�ϱ�
�c�S����nZ�c�Nh��9sT�D�غ�E��pJj*�gA0��OO�49��ߩ�w��i�Й������5�dz� �=�NGze���f!�����Q�k������������-4mG>v�R���qD��黥��]\������nG�`����e�+Va���^�	�j1��Na�T������#�, ��TV���a]-���@�a�}{��7�5ȳ��� 5 �oL�1���z˽��^���eQ�ŐT�w���Fem��|�ZO4��ÇWV%/7�R&�	�khh �FLT��.�$����:����2�+� {9��zpM�dLqW�3�Gvt��c�Cl�}q�R�du,Џ4^���|j�5�Q��X'��g�HZ>	Q���ή�_uH��#�M���n>�0�(Sz�M~0���j��Y��P��<ŉB.��~����U��=3��}��<�pv��+μ�R��<��1MN�R�]=S{��EX��1x_���R\{�[eǌ���yL��<M,؊��P�5�z�H�	�m�E��rO��$2���js���2ܰ�0\,O��q���1��ܮ��������r�K�������:�+�W/�?�WW�`0nh/��E�F#�MJ�[ڷ�Z�;��t!r�W/jg�rqvb9#&�A�}��W���o]9��6Ab�,Kw���km��rrV�m�y�hf_E���ȉr����Ğ�����I��,�}��1J$l���Y���o?�-�������m�����a�6h��\�]�l�� 1��թ΢H��mU�������?��/�o���MRr/�b�X�m��;m\�y��^����>'�}>�#.�<��P ΧzlD!!��f��Ȼ�3�6au��HP,��:���sA?;C���(�;(>jx[2+�y�n�~���ѐ�*��+(�L���^�E$m�Qx�5α깧�R�/e3��[���m5Ǖ<դ�Uᴂ�^!�u�e0	(��G.����J��|�D�}�5r�ig��.bѴ�7/tҴnu��QB(�ڜ����p��o}-H�y�(<'�)�.1x��6Mv�)�޹Ug�k�e_��s�(�s]m�G� t�K�+�K���R���/��4��UiQ<�g�^����{b�a䔄���;+�6M��x�~ơ�=�x�}��,��,����;Xv�c�wr%��I�E}1F��ȲU�[se��>-'�����tY���흛m���������|�ͷ]���&����QK�ȴ9�C��<t���|76H5/5{נ����6��saZ���99X�V���ǘ�e�[`|�CY�tag1-c�mL�~
���|-�����.������ɩ��͇YJ�ta�!�
b�v��vنs��G�uE��|�;��/�&�ԝ�\on���Y酝j��۱Wk�]�]�%l���.��v�7x��B؂��W��r��k��<ى���+���Q������iՙ�Xv��L�	�Mۭi�zQ�S@~�[͜3�-](�Հ/�|7��N+��\%��ٞ
ެ]�8����K	j���6\�b����W�S�hVP4�o��Rl��b�ȷ%&h�%�ViD�iR�~���@��&��=D�}�}A]l5���VO{l�G�n'[гT a��Ŝ<&�e*�"�IC. ��TR��^�M@�=m�b�fA���j��v�-:�8���?���p2J���\���"7ps�e����Xn|�#,;���Js`��t�L�jF%��{�@6�̮� ���䐛��j��"M0SC��莳YE�Tg�4���N�.Hi	1�B.T�bI�����؆�p���vg��J��Ό�PE�/� ��R�-U�m�6Z�m��m`GB+�5���B߉4
'�l�p<_��v@Y��,7����/N��{��7�j��.(�k2��Ȟ�'��}E�w�g�|�ϥ�U�J��#�`Z����z�.���ݫ�'�5��zT����Yw��á����w)�|�oBC|�����K(��/�-CR�2[����������R�h���2�cQʠB��Jd����������=F�bvp������j"y����d���*|���lmU �N�ۣ�����ׯJ�N����ő�7l�!�ב e�g)�)D�n/�!�J��䛮�?y`/��S䖀��Ö�Z?��^���h�S��9��lb��v�����x���H;��k���3� ��`tr.S�׵rB6�m>��J�G%��H��TpH�0�����,t0��%��������u�����Ň) B �p��5<�ۥj;���!�b'!\agbazx���]��\D�zj��{<ǇpǗwI�N�oM=ݰ��Zya��/ª�ޠ�~^����sh$Q(d�+P�řr�I���[=z׏
Sj�]lPh�m��ױ�Ǭ�Qڧ�L:U��,�8[�n7y��_d[�`�X{.ޏ�^��o(u�o�`�fQ�,�&A�Qn&�=NZ�f*�.�u�$.�}aϖ� J���2�\K/rg�%E�}:�X�S�jU��/���;e.�}}�m������6r�#ee���}S�~j}�s�mwJ�=���nx1f���B��ڋG�e���N�ю�}�^�-%���:�˟��~�!���>��&�,a ~>���f��F�+������.sZ��'���v�^h0�e��0T�6�������O��� I5J��|}`p.U��jb��≵���[P��� dk�b���R9�c������.7���v������$$���|__�^�;��
@�"WVN�$w�*�_��fu���!��t�|O�y�Zp��:EԆ�"���j�:�����go��"����\���Td��I�=���������)�-%�/_�����+앒���g�� �8_]Zq��7�k��]�fyR�C��nL���k���]�־�I#��J���y 1��s�Vc��2g��lJ&�����fS�2�h��E�a�4Y���>�dD�-�dec�G9V��L|~���f9�jTdO�'qlP,dse۝U����_��3�[S�@������ ���CP��*��K;z
���W����{����{��]ȝ}Pt��ڂU����ƀ�a��C�d(n�*�Ff︷��v1���}��%�0=�ߦb�#U��"�Z 3K�}��Q�*O�;�����r�2�XYY�dd������Ϭ0p�=K�μӗh>� �m����ykX�V.���^|W��wª�B@�7J����L��b�6��P�3�ϊ�(h�iɁ)����>SiZ5���y(bh+ƀ���M� �A��d7���lz�X�>��rn&��ۀ-(�BH�ٻ[߼��(n�������	0iX�d����[|N�Btŭh��������wte�9�=:J�і����X�%���R�����+�O����Ys�$���| ��~fO����l�M':-�_��=6�)/����ּ_C4@���C����^Ԕ?��ػ%�S��8z�#���x{k���-��1�3�,�gz@��5?���z���髠�`��L�ЁUĶ�?�zH��j��֌���㡊{���[ʟ�ź����F�ܔ�Z�- P9�(Ѩ�3�qZ�o޷ƓK5���(�����V/�DM�;V��IY ��7�G��`�o�M�v�2t���>@�{c��k� ��ŭ���t1�ij�s�N+b��bN�����o��N�
kf�$�b��uP�0�q���d��&ec��������ȴ����:��7w�Q�P���
aP�.G�k~^��/��d5����mC��
��YLLv���R,�^�T�E���z��O�1fAbª�\��_�RY ��2sL��#�6�l=��S���I��+	�"J�XJ�ӝ�����eW���g�(����/���=�X�3,7��ڴ��5l�ak���T]i�po#5��-z�Y"�ˍ=<�u��;��فv$�{"��w���\���Q�P�ٰ��- �M8�c��j�]6���2��~,��1�һ��ͺ���h"Z�W�����.£	'�f��G��Ɂ������~�>@Y,�f����M=�<��?��Z��� �_��0%�"Hx!��9Mo&؉���~�	&nU*������ZTL�x��^���� �ǪfaS�G
_q�!��;��\��f�z�ƯX���&�j�ݿ7�	���
�J�"�������Ku7��������	�x�N|���S!��G����/3C//�����U�O �k����sb�7��OY{ ����;�ϓz�:>�T����GS�!{Yhk*or�]��վѺ0\��y�(ۻ��(_V��F��M�G���C�����LOB�mA���:a�(�V�?��Ò�e?n�z��)!zpʬ�����}�.��C�#Xŀ*�x4�-3&y�����FB�~��gf
w���ͷ��z؍3I�B�c�!w(�k��yϞ�~ u��UE�@w����_k����;r��acph��9(C��ޏ;�76Ԥ�����C��-�33"vF
|k�q�'/͍�{��o�ʣ��`�e���I�dL����a=������A�Jȝ�����qRU0�"}uu��y!�sur��`b����*]H�R#���\c��I66�H�[��#_ۏ8�9,Ou.���鳀@�4p]𖃮ށL��=۠0��s���_��(����K����y�%i�C�2��7���В��׷���,��V�A!��W,���@��t�`s9����%n	 �3��T�D�)O�1L���7��E�?����,��{��$~�7M��6E�d	��ρ��^�����3���ȵ������I�B��0̣"�X�B\���䍍jt��$t��`�7`0Py]Z���H���QȍD�P��c��V5��WH�g�Z#O1�&2���|X�CG�RM��nJn
�#�_����x���>�v��xA��1���ѽ?`��Yy�t��F$_��B]t�UI_Y:�f#w_X���5�m�䏸RU���@)=S���N�I��T8_f�wWb>�HL��j�[��*��A�B�y@�,m=8K#r6F��E' S�V:�3�q�i�|�'���������j,:� n^C�� hF�.M3�}D>���]/S����e صeCB�2H��i'I�z?������6i��Ρc�:}!���ΡS��'��HIEI��F4f�Y/�5�YO�2؊U�x�DH�U���/�s�lG�K�Y�w�1���,U��&�Ӱ��S���#����xz���D�sv���**T½��-c�?��Y	@�DjS���1�a���`�
�&J���8�z�����[��G-��� _���k���d�iG�5�\���K׎"cY�]!�� I�S�U,
�h�C��ȃf�7���k!T|� �3��;�����Њ��v�j��������R�����h�-G���=!G��@�d�1ѵ�g�mNx311���޸�>Z�:zT��:�]�ȋ6-�h$��cx�&����N�h棟����r�-DR�8VP��J�����$��S�P���Mo�M2ȅ@�G�P!9�!�&��DO3ð?������Lٞr��v�T�5�l�GK��nq���\ˢ���B�0K{P�0�9�wrt����h�=�,P�)kgUzj��-�@���c.�(�9�_j��E:��s���4�v�0����ֺ�X��Ø3�+��`Y�S��̿�F��u�=`���1���a�7��.}9��WC;�?n��V_٘+��l~������?!� �H���j)��q굡w�� C�gZ<\KN����������Ό��
/��ۏ%&-n���B��+M{�sӇR�o�@���1��[�<$t�1�5���=_l�~��n�W��Е#���6.�mb��[1��I~��b�~�ͨ쎾ZK���so�&�4�D�D�v׃�p�#����P<	�����~�'ha���O�͙�z���{�Nת�Z=�D�����ol�1˝�iW��]��MKFD� F�o��)��q����|�33l��M�u�a���)Ô]����7�d�f�����G>�h���Z������$�^T(Z &*����.�̷���N����ơ�
�b-��ߓ�v�O��Qd��b߭�^����Cn��@~���Ac����6>Q=�B�y+�MC۞������A���RK&�pS�K�g`:��#����#H���a+��Nt"�p�q�o<�܌�6��R�!I�n \.H6�vz��?��?V��OX�Q�`�6�'~�ޗ�0s_}�~f�c^�)U��0�y�@'��n�W�� ��I�OÍ|n�8��m]@�)�C�3�\-�F�4�gx�
1����Ί�Z�}������)�J@ȝˮ�ݫ�#-�[*��`���dɹDI+��`��Yb���]��Ք���nX>�PK   ���X��6�  S# /   images/ea543ea3-2b47-4327-947a-6d32920e175d.pngT�cpf�/�<�m۶��mۘضmkb;����۶�Μ�{�9���޵v��^ݻ���
r�p���@@@p�"J@@ V  `wH�?+�/��NJ�߀j~� I�����@����<Tx�O�:%��;(��RFFF"��*:�� "�*��'�������������ϰ�s���Y��{���=�t�vU��b��vU��u�L����%���BЃ���,��3%���KIq���Y�d���!��r����
�������?b1�ˈ�/-� M��AMA�C�K��Ƈ�/w���H[����^ l�������1�oN��2>���_n���{�2e?�3Q�������������6m&����9��������,�'������������"�.�^lM5õB.׾��+���:7�Z�<��s��Y�dƱf�έ�\(�KC�հ(�v�őh|7{
k��R2\�����T%E��e�8'��B��A�����=̩�Gi��뜣�f��eE����V�K��J�WU� KК�ay���__ώ�)k�cP{����؜���S톘<�c�f������.x9�����F#�,��t��_��ʭj]�����r��Nk�<�i��bɔU���Sߐ��p1raH5�Y���C@��Ӡ�w���xz)�[kQ�5�Jr�SM��w�lMF�'��)�M�˓���n���s��R��ݲ�Z<n��;#D�f�.�{�>kJ�ny�%���c!a�հ��Ģ8��G�u��bB��e�{��|�͵�P�G���=I���ߟ'��b���3��8��c���y��~�S�TxB���%I0�ŸS�J�i�<Q$ i�%�,w@jg97�4��7�P�i��uk�R�N+t�I9�?�$���|�|���
 
Ɏ[�eBJ�C�Ľ���G
?�V��\��1��5*�f^�r0��"�x`[��s�f#w�����o���Â٢�I��9��W�&y��B��&ր[Z�ở`�+r��	�D��M�M7�e�8œ�	|���d���D�w?m<? ;��=�Bf{���>&��w���*\���GO0��$���K ����8�'� \k����&�h�M�#�3��	\=7lN B���V	%y����BW�Q�pu���w�A<M��2qĝ{.,�f:06"�+j�JdM���1��ڿ�bJ	���`��3h�5��`F�¬bE��f5PBx�8R����M���"�I�� j�h�+m��A:%4��M��9R?T緉A����U�D�������pA7����c��m�@���V�kp�H3�7d�GQ��D�:�t�(�̈- v5�	)G�Pr�7	b�[^f3�x��B�~�R�7c��^(�lԖB�dB 2�D1�~�5��@Ne�HK���m=x�t��&S���]_e�� ��J%@�Ư4Z���0Jb�(R���H��QN.����ް�`�4TE�^8�w�Q��	)U�!$k�z	ޟ�ӳ
ku ��r�j��Vz��iq%�/�G�8�H2��(�A�|�^t/ߓ<���T3�|�r%;+�Dj-Y�<�4�ql{?�(����U�ڦ��)�?U�n*���{�V�9m8��҄Z�T�CѨOJ,9�F
�L�X3���X@N���`��-qDԊ'�;�@	`$� ����fa�mE���A�F6���PR���LN���ɍ��{W�$&�&��V0'��SX&�������y)�r�JF� %eO��G'صމl- �����/f��|6����W(/p�
!���3�4Y����~z� �w#6^�[�4ɯbu�S��b�!��?Ԩ�����q�K$hqZL�D)O�x5b�<���G��^j��!
�v�'Z��4�cu�7����_�u,�^S���v؉�&�x�AU@�={���6[����%ޱ!ֆLxZ�PQ&�!�3��#رr��X�	��BJ�*5N���$�O�� J佄R1"Ղ�������c�x��T�T>�K����9��l�_4=;],X�-���܀��]tƚ��[GĤz4�_G@p��0_K��?�p������o�����k����o8���Ө��yyпr܈��r��s]���{?�!@&2
e��'K/�!�+��-�%J��ycl�᠇���E95k��΃�%�
:�1@h@y@Qw
b��g/��y�|d���P���"A�R��_PGÛ��6�f�k�P��TFN�8�nnb���ϋP���0�]�V3�-��K���7�t3��H�8�ް���+D{m��1��Z�L||tG��o�k�+�Go�Hc/f%��cb�\�jN� ��5a���LL�x{"I��Ț�q�}���*���px��n�o��> L�����-u����W���A�_w1��3f�IvB��~J�r]�� ��YhѴ�5�m��V��GŊ2hM�46L��nH�D����@q4� �m��#ִگ�Rݕ�5D��kP8� 0�ҽ�8��l���L�e��9�_�aZ��ȭ�!�Ķ�(Ɵ��'(q��O}�oW`�V�j�;=~�5���M��ߝf�ͮ������ٺ�4FfŻ`@��Z�#�<� W�kB�g)^�ްq���NGvq��BiQ���S%�-�o��� ���z�-X���e�I)*��m���t���>O ��QEc�� ��9�z�*�"J�7����`u��$E�Nx�:^,�Jo[.����u��2w��Q����Ω�<����g
Y<'�����?9`����3���:H\Mgk;_�*M*o��'vC]Ty��/T��X"W82�2+(�"�(���fA���`a=x�U=M˚+Q�Ch��b[b�X6"�7����!���n�*���F�j����W��Wt 8W
��"�n��)KX�T�3(=�^=Γ��Mp|w��@>'$|w��G�l��pHP(,\g��Wy�	����7����|?T�g��Sӵ�.�	#�v�ߛ���$�B#�z������Z��W/(�VZ�B�6����C����Yq��	���l��+�uJ��5�%)t��k�8����}�&X:jѦT�%��J��J��h��K�?���e�u�}آ�ubt[t�����LqF�����_ې�7~�+�6�jq?)���@4�C�L)=�����9	�P��W�m��'�'���|Տ�_�gB��$�������a?��箖����E��!���m �}�c���f���<������!���b�`��_�x���D���g��@���s�����>�N�������=P��;�N�}�W�v�/�����'����Q$1���>��nn���Hp�an� z�6;6��B,�OO�n����)�R��ܑ��[ӌgw�?�0h�w��
�,��%y���#��NRZ�w���V��������$�O7����l9�>\�by�&3�a|��c!3��%I��m��������AE� ��\8�yQr,bN��0bA�[�cLW/�DN�����tLo%���Ե�]�Tʄ�6�uX~v��`�d!2�j�����bb$�ƻ��w v����V��w/����4V�`~5eS{C�x�`e���r�t�aD������z����X�j_��Q�[���[���\��e�Z���d���-����O�+�n������o�C"iO"���:�;c��ʿ� qU��5����aB}t\v,1�˒��8_�+��I�o���]WB0q��d�J��'7�Pd���{���}~w���m���a`��)J���4~$G���������B��xc]v�3v�5B�
�@f%ɽ���2��QD��OB�>ZC�%�����r0*��\�
��� S �H�F�Ӌ/gw~�����i����O�A�?���z尻{;:Ox���یW��I���K��vQ��@����626A�����~�������7$%��fBn� � ]�����b;�����n�A�����r�g��7�_H�C��BV [���V~�𳠉��/P)�Ex��^�������u���������S�0~
���sW��d�f�K�Յsײ	��Wi��rd��aʲ1���؛{��T7P����,��1����M�O�~��X���W��󻳺z��=�'R�>�*����NC$�so������ �uz0����V��_R�� Ԡd�q��;mpA΃�m<��8��s���8㔼�Ț���Cak��-���_ԑ�*.e��R�v���@Ni���7�Z����#�z����빞!�w�	����?=x8�}����)�Ș�˨�^�k,̎�"In#��en�DibA�g�ɣO�PH��Q�a�e�j{5K{p�zv=ұ�����; �L�΀(r^���"Y��p}?�������s\x�{��L�8w��gc����W"��Ш<r�!����F�b8zv�5^G�:������@-��o��i���������������~��&�����Ϳ]��tG�l~�;�#�q�)k���pf��w\D>�~�s�BQ�}:�^��AJ��H���*�]���D��O�l�ӹ���}�t��ڄ]��.�PD,\��zX�mzM��t��w)�D1�Ak�u�����8�4c�m ;TUd�f]��K4�P7Z[2%��?���K�t�yA0bN�T�_��Q�M%r\�,ي�<��T�|�����ݦ��p���Ķ�+��!�ޟRRv�H�f�i�z�XH7���S�$�ɰ����Zc�8��w�_��@)L,5bsL��+I��-^d��yua�����f�a�Y4z����ANfi����&�����i�"���K��ZT۸^��f��������%�J�^g+��L��հ�>dm�#Ͽo�����o㧂]��yB�W��g������΢W4E�+�I�}}o�A�^�N���c��.��v�P�<]��cl�N�Ӯr�3��j���Wh��Lj-��c�I\U�
��#-0E����ʫTz�FD��;Ʀ�6������|��u_J����K{���/"���2e���d#�f����'is�TU!��I�d-�Z��N�>⽇�&~�Y�����fG�3\n�4�g�����H���4�����Z:�{���J��ր����i�YZe��� tS��qm2�O�д^Q	��u*u6��ұ����8�C�tF���,Y�ع��!�/���SΗ`7�%s��ֵ^ASD̂5��=Й��1�C^q|`�i��k����������nq�E�h��3���	�/��f�F������X���� �K��+�Z������^ѻ��9�_���S�a{��o��o8�Gp�yk���:�ݾ��0u�������1\�ƢeA��>}g7�wJ��$;G���Z�`�ۆ�1���j��a88d�8��1���(�(�~D�49.�h��C37������3�]��P��\�� w�`� D�Bi,YrS��>��fLuJ�G�S��ƺJ�]��td��(�[}���1Ov�vs��<i�74Ɍ��S�Ȁ>r=T�
�h����jM���.D�E�R��o\@��	�A��ы���4������$��
S�i�Q�0N2�H�P�i����ioދYf����<�\�����d�����I��$
�l��[���%�8N e���bYX�/��Y����7������8j��gj�;�^�Z7w���kŝ�~�����b���;��oz�1�/�Q[ ��;���=Wə��C��f)~@"L�+p��@8�]�$�2��Vte�'���!�^B�&%W�CT��;�e瞫��g��@�^�+� N,/�Cz�Oak>;�%=Olp�u�/�?��<#�9��cҭ�>�i
e\����ū8<0�1�O��顇O9�q���vJJ�c[h�K���޲e�K��Rڧ�Y6W�߻\���ݡI�3��6���j�t��d���JA�bpI"U�H[�����&:2>�U2��F���s��$0�`��hE����氉����{��^�Ι�º��P�mn�g���&��y�>�e�O�?������,�BC��5{ڗj�v����P/��ӕ8�#��9k�Pr�XwY�"�?M���n�^��t�t���X4�<�����f�=�v�-�m*=R�	ʜ:��~���2)����Ϫ:����c��������5\:��<#7���@4g����cXG��<t����L�0y�|�D��z�u��@�
�����7׉}��T]�^u������X������/.��\$�J1��D5�I��M��jN�JF�g�}r��VH���tD�ߖ��PM>�V; ���E����򘹚_���Y�C	(��~Ph�~=x��w�S`�.��-��6�S[���b��(@�`!�!Ô%��ιI>#�Ѹ`;�K���$\�fim击�-��ﲞ����n�����Ng�c���(�|l��yv��
� U��N3��	f	EڴkI�Sc����*p+�;/��K]�!�}m��������ȕK1Db�9����7��n���#��[ntz��6�����򽏑�W��5�$~��%�41�U��G�󶣞���P1c��Ȩ��֓��ۉ�`��~��&S�����kx*V ��8�e���mS�:��L�^����pK�'�->������w�D���CW{,K[�6n�������{�W�9�ܖt1MI��2F8S�"s�Ag<��Rl7-�cf=`����oę��.��ʻo(�NM�����%��'*7$�F��C�ܞ{�=vt�cXwXl��l�Q
�8};f�	�̯�@cf�K��"�I��3Kv���du�4oʽ�.[4GGGK�[1s��F2ZO�;�x�����Y�|�Sߌ�|�����{�}����朅��x�'�����ji;��^����Z��D��d�c���l��ia�m�:�'��k�g��"(���Z�fĭ�#O��c�̥��lF@c������*��ޝ���4ϛ	�� Ӳl�<_掎=?q=&�� 9�˻�s��ҿQ�HNR�V���6<���~Z ��u����z�a�
����6t���q?o�3�}}&��<��T�=B"U�*��_�&u|�K�c��EU*C=�5����]W��s��z)PQ���)���*���ٌF�-��w=����<O蒬���-A����� ?c�M�O�X��Y
~�MbZ�6�+o����2���Z}nI��8�ޛci&}���+��ų9c��z�\�%3�&��n1�����\�mL�����=;I�!|;@�� �Ĳ�n�u�o+���$&6k�a�T���}>�B����hHЄ�f<H1����P��!x��M��J*j����B�Xw�@�\�WN��n�u�gJ^at�\T�y�_4���|iQfҝ��`k�� �h���xg�<�X�}C����h�g屹G�����ּ��z�zlb�lJ��Ilm��Hp����wH�Z4�_"���۴��C���G�u�`-$�Xɕ��pN���N�$C�MS��=��)����4�Fo2	-�~y�w���d�'����tB�㪧��\����.��p�ߎ����v/��׍1�\�٢���ز� iƁ���N���r%4�9[�r��Є��gl�h96�Aʒ�M����c�*V<T��&�Lr�����$3�"��R�/'q�H�A]t^�j�R:Nx5����N�Ns�I4ts�ş�ҳV��gt����X0�vl����m	<S��тVQ�τ�� 3�$9�]�'�T�����R{��-۴�\�*4�PL����q��n;Hm���Y
W����1ouܲ!U�Kez� ���)�gP��ڲ��(p�Ѻh�tS�[��>�t�K�/�Չ7+%Y�+9�)&��� ��d�f�/�c�7>��Derl��b�e�F����t��u����kƺ���!X�꼼�~~�4���K_��9fv�vw��X o�_�Y��sY�«��V�ax�!�-3p(Bh�Q����K��c��&���Y���qy�5T3Z�J���$\`@(�`�2�\�������D��D���F�<N��/b�#��p&^��Tį��nӾr�b�nں�����0��B&����[�F�#�i�ҙ����ȩ��aq�����/x8�J)��e�"�3�k���LԤ��X3�\��e�B��w��Wʸ�"�]�R�Tu��b,��NcBWL�'�;R��2&���B��X�.\s�0������>(����td�e��\>o6�e��@x}��XD����谆r�4�Ԯ�y������<4�����z1|��.j�'��blo� �UZ���D���)��[;�0��~0ᠰG����`JtH���zB�01���O�bA\D��p)�qB���Č8��G�h�]�)G6Y}� �:�UԹ^��|PN������S嗩�W�k��:Nd�RqI�^V���6��b��(5'�F0����ܹ�$x�����M�WLItz�1i�����n�Wr��TIQ� wZ:l"+N�(#U��(ۻ�Zp�b�F��H{����f�[�D��b�2����7Ύ"u_�����:3��Vt�Å�L8��[��0Bl���ȺeL@IS���Ӵ�N�M
-�� ��5�y�������G,��o�d4O�/2�����^}�����n�vd�h4�ʚ,�N�/�^���D��Ӓlx648af�6'��_�S,�4��y�DJ��=c�^|d��&����K����F�$��2-�Q���IG�=�J:�u��`��X�A�G�������i 5-���F��Ϩy�zfo9aa~���T��L�)/���$*[�
�9� ��GuЁ��˂P�QTp��;|�*��r7��D[Z�Z6?QIf��C9�䰎z̥7�J����V[j&?�V�9;z��,�9m���?w�Dq컝ix�ܘ(ǅ��;�"2q�,|�T'������M�;Q��3��������?1�O5�{ۗ�ںKz��k�ǬuC
��VF���B@3�8H�F�C�SƅZ�Ȍ�Ґ�(�;QȪ'���S�%KuN*�h�P����m�-F��K�W��t��U@"?����͉�9�k �����IWy��0�$��������F픰�K:��ɍ
U�U?�
I�� �O�?�y:5|�Ht��-�P�{*d2ڼ��^��;kُyC�/��C誂&1\jo�"���u݌&Q����h8���:����+�������\��\�rT7�מ����%�T��WiR��dWXmL�IZ����ÿ�˃�B��Ճ'�L�6��߾���.��}�u��=����fG����O���T�ɀ~FBv�	/e�m	8|V3j�v����%�	�K�QM��b�1Z�"[�I"U�񑒑vE�:�a+��	O
��fS)�D㳚H-�	e;�+j7
�,�����	q�Pԕ9 7$sc^J2ad18���K��!���� ���-+	���FG�oG�a��Ko/��r�[���V�5["҈91���L��¶�b��x�E��<��\IU���0��R�N7���?�����|QB�	��2�;-YZ�	[8FMfd3�9&�$Ou�V"���d����qT�Wy���ÙbD��	�#*� /�P������`my��6CA	���e�����>1��s�|;F&�nT�)�5&� +h�� �
|"�Jnd�v�d�֣0��XT����� �=ҁ(�'�w���K���_32\�>��,�����F�Ut�`�_��M���G�]JBL*x�^�L�1!4���`7cF!vM�6��&<=-�/��`|^;��> PJ܁��H�~� � ���J��VL'��7A=V���������BFf�yF����'�p#�.�Jo�k.U2���G2$�� 'p��}Jů4џ���H��?Ԓ��:D������j�bz�f�fCv0\�f�L	��E��%�
�J���>S��ރ��sk+���of����~el����/�s�#���|��4�ENAa�Ⱥ�s��9~��A��(JA�.��1%�C�r�TPI������</�,Y��]���_�(<'$S3EĒ��/��G��Z����0k��:�x(��L���/$�K<	Xc��2� �������P��_��@�k~�Z RR
�!�FNtJ%�7�bB��B�;
�ꠥ0���6�=�(��ãϑ�k�gU�GQNi"�D�2��'#�rdЕ���%�Yr�4�%�#Y��o����N�IQЕjx�ʒ��-[�X�mפ->�W�f�	dT��čN�aLص\��y��֬���# [�S��m/�������}�R:�4�]ѫ�b��Ș�cm�ԺS��~°���ѣ��%Ե8����Dm��v�R�QB�s
�X���"��c|��ZP��ZE�x��\8���\IF���@�n\��6�l�WU+�遙���������ų�b��$?���+Uk�V�*I��숊�D��3�|�? 	X7J�A؟�߸��Q�x���9�$5IY�i�Xqn'`QT�M.��������5�k�~�(����&s�Ŧҝ�Sښ��hJmGȈ2bfC97��Q�9
U�M��lK;��v5M����;ѮS"(���h99��%9�U�&(}�KH2�AS�X-1� �y;`⋕�����^m��3\Q�`|�~Jš�?����6`���
���?kv�x�PI����<g񶺏h�m��P�c<��$n�$��XИ�L�g��y�N�6W`�Ǆ�\��oE#d�=������*��SV�]��RbC`�� ,��N��(Np�Bi5dH���	�m��9�hE�=��T$w<���eD�R�|KL��~�@�!�i̒�l�M�uĂE�{x�y&C�:_sܜ\�q$�EG�C��2Z}�[��%�$(|�9%�:��>�	���̑���6��&^
���P�QEؓ*�Ҿ>3���z�4`�K`�kk�b%(�e����U���e�T���&��P��4��Q�n����U?�w��,�w�?YÔ ��a:�h,�U��u�A>��F��(6��K(�=�O��M�(���ӆ�t
y�2��ȡ���T;t>z���z:�O2l�����X%���%��J|������V�́��z�Q{	�h�UF���f�{J�ZƅJʧ�C�U�@\�����5~���|3N���ԧ!�~4.ދ�v??5P�gGi��v�)eQ�365��H�iE0�S�}�����s�JĲSaj�mT�i�`��8���غ���YJ�mHYIHӡƯ����5�����Q������"a�$�f�_됸��Ci��ǹx�q'�Z95*�7�Y��K	":��
��`r��ɇ!0]s1��f6�3-Ǫ�@�m����rt��KZ������djͷ�"C���zV���_����~h�T�R�A�Q�h�?+��tYт-7�F������Zګܯ�2� Rv�Y�
��cۊ
��䦊@`���<r��4K�4�'��o@H�*I$�T���/ś���X�e=�t�h LK���|����DC��b��?w��E��NzI�3M���y�[��?�?B�� ���Jj�����+������,�s�6�`��r֨Iosu�0�gao88�γ(�QyS8�X�W��L>���H��>���)=)��6H'�y�3ߦY�y�E+4Ś�В�UE#�沊�#{�7�����S�����\�!&��l{O+��E�� +�mav)VZ�i�% Iu�)�(�g��-������ڳ��t�3L|��*�����{���dܺ��U@� �D�������$t�� �r�<b<���*�
�!K$*��?0ܼ,h't�C:֔��hZї
��ڀG,��S�G��K���y�͠1B�.D�v����1�!�1qݘ�_H�eb�@
���'�ӭ��a��W��Mm���RQ����`�XT���@����O'$b�q��b��X.n��3�M�f�]��LE.��
`�ɾAo�!��>īXT����E���%���CŃ���|�o�����P�ی�1�	JG{��~��'�L�G?��Ih�Sў������}��]��U���e3P*z��,n�������}ΖI��+���vtx�mݹ�$H��7oN�"Sꕭ��CkЪ�	)W�j��!�x�x����\
8�b����i�cqG��kw'Ӱ%���|Z� ����e�Z���=��ظS��eO�;;Ц#��u��9D@��Rc���w��: {6|�?Yw�f�Vn��G��1( �u�$"ܩA��l%�����Qo��69�����T�V�	x�)��!u�L��ۑ]�g�ʠ``H�˰��k�xa��'2�����ֳ�"`oa��K��$x���0Ň�"ȼ����\}:0����]Az�(:�3uQ}d;�p^�|l���d F�Kb=���GCrz�;.{-jBs���'+��^ �ݜm2���pq\�tW���L}��B����f�� d|N�،��d�e�Lc/������i�R�������q]����w@���=h,���Ǖ����f�C?��K������K�*���WN��B�)Ur�yWV�s�(|_9u�!�>(kbn��^hռD�0�j�U%�ڜ�]4�}E$)]��B=t������U.oq�2�zHŪ��h�"�J/1��Ѹ藤�Ȓ��2�Y�JHv������H�4d�ﺓ�L�H
��&y�5�g �]=zhj5^�����4����kȳ�kC5{��T��-��C�C��*�n��Vn<,�N�{�v�h��C�)&���pw��P"�p�U��St������;��j�:�6?�O���W�l��g���.����^�|��~�~�HåY�<se�灪"ğ�.;(�E���*�
�\\̶�3f�UrB_c4�r�ĵ�\So+Ʊ����o��c�T_�����
�R��}d��rqI�,���˫��
2Ц�ˆcP�*+�?fRT����3��r&=kz$�S 4`i${3�F�k�ޟD@*&M��Jx�����s�����S����-4�(&C��M0�p��+hC��$��R��x
 Y��-�V��gT��ɖ�d�N�*G�{��m�_%���H��W�	0�Q֠KcU�V.4~oƼt�~����
-��Xή��M���f�UC�|�f��[��ܭ��d;v5:�9����?�[��t����ia���T�ʺL�bD-�ތ�!t�_�Ầ�ˎzBM���gq@R�IL�y�_���qo�T%X)����~Wq��P��9�Q�i~��c��A0R�r߶�C��w$j@��$k�j��қ���h���J���t\H�!q�Bt�o&K�
�t��rrC��.A�vڑpU(E��PX*53��v�v�I6.Ѻa����)�`�����[KR�=�̯b"\��#G|W�QLE�>�E�KQ+��x������4����W��$6$���X7M��a>Ǳ���K��̩t^��n_�X٣)<(�e�,` !Ws����溨̍:b=f��Ԟ;qK+��$�_�۔y���sj\��������#*��zjH+�J��_��K��b�续��Sr���jTY��B���
�r�h��:�K���W�L��BK�>h}���s�����jthOl^<.���\WSEY֑d11��$��Ƒux��E9�ѭm�Q���.�>9/^�m�˓�  �H��1�1�\�-����r�u�	�ʺ�B�-|��}���w�Rn���,�]�̩����X?"�>��y�Ksl��u��3iS�N�h�4C��v�#;ǝُ"]CUp�m��Q�y�5R�i<a,mj���_��|RO`E��ʨ.'��o�&��q�]�X^�.(Om乚��;�@���ʔ9k)��u���O%��lpV_i�@���fR@l\ ,��T���{�gb�/���G�������m}��EM!�V3�<�0�>N���!��+�p�hϤ@y3�S>�d����$>�)��s��I��A4�$��Aε|�>�~]	J�v���\]���M:��=�q�0�c5;���#��hyۜg��b�~�]�B5�}����ui��k��/��^FM��Ve�&.1�g��Az�ZйS� ˬ�JG��|8�c�|V��4�Nǿ`�l��IÞ�E��6�_�n���4�\�ǁ��x�
_-Xtd�0T��k0�T���0�4��\��^jP:�9�JZ������HM_8�c(���h|���k&�ǋ�xE���^�wp�U���" ���U4�i���j��e-_'�LYL�*���`�
N��q���&�d�e)��(M�J�={c� EF뵔i���"��O�F#*��O���>�9�U=����>A@�m�a��r^�x�sJ���מ���ڊ���':5���ɜ����*�ArODM86�D�U'y�ƭ]�/�e1Za���6~��{�>�:s���^;��f$iW��D�	�&�򠤨\����`z7B��}u��X�'qbe&�Ĩq�iq��6��$�My���k��o����x>N����`(I�掏��b�ɺ�ݢ��ߘܧd=nQ�Ĳ���]�-3@4Rh�ͨ��~�D���;�q#	܀<�=hO9
-�,�72A�*�?�J�Z���3G$3t�'I2	4h�iG�,� &��N�����k��ч����&O�' ���6���Э_`��a��)'��Lp]�uYK��2�~��ԉ�N�.y/��f��GC��?��[���)�¬��v��s�)�n��Hg� c�
.EjW��u��xH�PYhROj�@�~��mt�&_Y��{��O뵂\��f��b�oP��2Ա�8~q:�K�+&��*+��$ٜ�9x��ѐ)O}o>D5J���Rrʳ�K�E>vrs��&'��8�5���GG6G:UyV�.���cʽ#oHv�L���5�<�S�0Ԧ;�n�aeR���I�����^|��N������LR>�"���8��ƞf��b�Zj�t��ֲ��5�H\�Y�#�����jr���P��aRkV�z���jn�K�C�PՀ3�d����`����z��ozKB��� Vl�������hJVs��~��r�E ŗ��Eǜ��]�P�&ng
�ڤRV�f��,���^?&�C�!�4@�v׳����D@0�z#�S>��~�Q�2�	w�l[<��k,8�fʹ����ٮ-����K� X:
*)��m{Y�{ 0K.�(0���j+P����_����ƣ�%S�lvU�q�;�l�c@�#�΁{N4�>0�hB�\����`��n��+�\�ޤ�Zuk|�Ba��0���y2���fs�R{-]x�l�N�� ��t"�2!qbY
C��a�����-�.�{*k�W��&܂�l��Q��e�3U`���c�ŀ�����F�'a}�n��#�c̅����1'*�t�n��>�Gl$}V���7��H����xfҿ��MAX���i��!=����[cQuHe���y�_��
V�:N���'��Fqz2�2�x��喚;��x�
֒�[����ѡ�x���nV��(&$?Nli:�Z�I}9*��L�\G��U��$ȃ�I�q9"��X�IS`D4hъ�"B�E��u�)�����g/�wm�����X�^3� ���5�m7�jn�/M�-J�S�e5�����Tg�E�x��S	S�:CS�L�ߪ��6���"V�EoL8�.��<SĖ�eW�P��ʼ]�����T�*��FX04ڷb�U.P�*�v�� H�─)DQ�lEƪ{t���� �>�nuZ��yySuU�ᓹ�Ԧ*2h�C7S�v��������zؕ�Ηq���,a�5<��!�����zp8�C�*�����=%��̅�f(�?X �s�`B 7�hD�������<bw�s�C�R$�|�@������F�]f��|jZ�K1���DU*Ug.��xR�N܁i��I-
������l��n�y]��Fz�tl|n�J����Y�A�;:ڞ�z^==�M��9!P��LR�<���W,)D��~�}������<XI%q'&o4[�]�JQ75)��� �ɷg�R>@yE��X���R�y0�+3��7z*;�����{e�up�<NP�@
�`��߼6�	�E���(7g��P�A,�
9�J"��o�G��jǧ8@K�`��db̄=�N�� E����b������B�l����VQ�(Ƚ�dY���sy�73���yx�g��2��.{��8���Еt �&�T��}F[��AR�/��o�B�Eg���y���˧��ݳ1�M�k�6#�z+`_�Q�J�KS/"�1�b�4�c%\��۶vlg�6&v2�5�m۶mۘ�6�{�����UOw��w;g�Ft����H��r<`T��$2+Q>�E������ߧ�2����y�<�`,�`
#!�!4AH	E��kMuEC� ��͜ea3I�yiX%p��
�Жl������|.$'�І������FҾi���#�f����86��_�ѻ�.1f͘>��"@LD���Z��LD?hy�fV�>��8�3�H�6��H�U�C��e3���r��_%2�NBdr5^�`��Gj6<���Lp�Ѽ�7P�ͬ�ϩ�A���:b��*@��K�nj��/.�d��������q�.i���=X����a��bɭ�X�q7��x�C�;��2�3a���c�T���x�ڎ��F,�0$���,$�+���RQ���F��\#T۫�����L]f��L'�;�h���Q'041��d���{d	LZTŹ�W����%��˼�Ǻ�ϒl�2p���a4�&�m�μ{��@�9t�	L3�I�Ϫ�<��4D@����%:��z����o���뮷�O:y�
��Q�iNx����_�Ҡ=�٪��Db�`�E�SWF[�^�k����5�H�<G�]�n��gv���%���~�R���Y@������+Ne�c�����.��z�Y�������N��8��5]�{k�.}J�(?Rg>�_4 �b���yUVr=^Ǧ�z�:Y�ȳ�ړ��㊃oT|#ZR%kLA��rFu����<NJ�2��۩��Ф���)���-
�2�]H��J�!�_�l�s���R,��乿zv��C�	[őe�f!��7���A�H���<�-��q�8^,xCSP�<����8�T�\xPï����Pf��{B���K�/�s��(Z���E-�>m�w��l`R�&R��QWM#z1�Q]wbDFR8�55�9ν]f�F�U�Q�+_h�n@�������G�J�L�N�f/$�g��f���$�K�����U��W�4��q�pp��o��l>k��Ϋ�d����gsq��k��l�����:�^���|�L�f,��ѕ��"_�be�C~��)D���=LP0�C$擔���5*��&��H��/�:?�:ya�v����W���eKur�II0��n�<Nd��C)9H_]���q�锶������1�G�Ĩ�?�)CH����[��(�H���Zڎ�K,��=,�s��e���e���N �~L`TƮfଠp� �"��N����_��
���i`֐<聤w�EY�[%�٪�g��3Y��,.s+!Q��K����J��S�<l�b��Zx���U��az��F�n\3P#^����z8��	p�	
���q�S��`��g��C7�a{����ݢo�����=!�WB`���2����i~�}�YNW��!a�}�%]�j{��%c���.����Zi��R	Q�r�%5�`Z�CE��E�2}�t�e�	o�d�Ny�'/���P*V���N��d��Қ�Q�Ӂ�>c�s��SK��"
գ���ͳ������T��/��t*pJ\b۰�ybs����x��������Q�wt�3��a�/�iyݩe�ڊlG!Q�>�*z mI�/\ޡ�/q�z�
�AV��b���2�E��!��#�</�SL=9om�B9���TV����p�@�}b!�� -�6�l�B���-��N뤴�z�d�00Aѹ�ٟ�T>��qy���]�w=4�����~���T���e��q}�G �.��=h�`'~וL=X�[�MW3��$�M�����@KkN�c7����BKgtu��W��8rv*A����dC�#�bMl�k�Q��^��cR]<]oC�S�@��v�	�f���i<h�g���+�D�r{� I����������C�_���tWH>�A8a�`Cm��"m$�A�mn�rg���@��lDъaR���
Ja���+�6)R�r�y��^'�ދ��C6���Bp�9J��	��,��=��� h���4C��Hs��Qr9�[�;�phS�e����\m�h�BlN=�p�D)���R���I�N���O������,��tqT�!<2��G��h��0/@{��\���� ���2������~0�y�:w��,́ ������	� c����]z-����(�J��p2g��`�[�܈=���]j��N&-,�t��ؚr��"?gԐ;���x�BEK5>LvC
�f��uLe���p��[��t͚N�M�<�ԯ�vrl�-�CƄ���|���kl��A��D,�i���2�#k�:��kSP%J-:3w�� KU$TѵA��+p
9�#h8֗�DsHͣ����`���st�{9��AwB�u�W��1�O�R���,�i��9����tE*�%���m��lAY��/$Q��.�/0Ui��up��	�)G"0
�*6Y�I�g�Ĺԅ$��D�1�r��3�$��{�����������;{#����������f�"��2��M�5����(�Lp�f��+�|R�����ӹ8 *�q�S�{�C��}	;`�����H��gj?;'ص��`3]K�]�"��ف3%��Y��OL:�����TsL�.���9�-]uF�=�,��Ԋި�W���~Z+`�f9�K��>Ǌus��ԫ��&0��J����%�Q�������L�U�@�I��X:� ��F_gx4*�Ū}��1N�p;n���k$));DO'��Vk�KĈ ��t�?�.5��lԢÝ�cNuC�#�ҽ�[DL&ck��s�D�>N��.Mh@���8���Z3!.F�S�r3X���G��}/w��yK����1�C�=�1N	+euh�]D�7}z�8(�U��l���OY5rvV=.���'5�(Ѕ��jU�x
�Q�j����� �Y�5��B�l�{��)s���0���s�����|+<�\��j�7��'���;~)�ᅜ6eTx��cO��7U�P�����0�S��3�"�4���������,������!!��&M�䓀�7%�Ě6#XvQo�8�7̤�Eܭ���-�߄W=�W�銤�����pV}�LW]ĳ�7��wH�n2���mPՁR������\�DDP�Y��|��L�i���(�/�*+`�t=1��7�6
�>���5.7�p�+��VY�������/���1$I ���b�V�E����f�$��o��`zRQ���Z�?޴]8���\�g��y8y�}j-�$#�d״Z�:��x势" �������� �Q�E�d�-���X�������1n��QZ��]L�/�]� ��Q����ܪ,���J� �ƹ���IV|a���F�1!�`�H	�G�?ˍ��y���^��ʚރ��j7onZ��AFm44lU�Rf�a��E��_�S�lJ0@9��_������X4���;S��x�Ё��>[R���X��"�c�T�b�m�Q��|A�D?�v�ͳ��#<E�V�"�:����>t���.� @A��N�P��s�5|K)�t>B�ǹ�(F���d��X��[�D�Ċ������D�fn�I��ѳ�>}t���C��$�c.V��j�"�I8ʳd�=�L����)���������N=E^=�2�_���.8m9�>�h<���(�5�۽�B�ѝ��4�WB�3�˯��H�7|_���oL�`�+m��:ڼ]wY~���2����v�W�G��2Y_F�h�>lu���&�OI{QZf�~�P7{@��DPr�ضX'4�^���5+�p#�����(���,�H��H�@H�]sd���ܬ�@6�������Y�d��xnDݟ��x���Fިbڰ%�1�*>������ �P�s>�E@D��i-'��+�J�C�@m-�׵䍛b.��c�a�Iv�E�,�E���g�=����ld�dx��O�(;�9��1T�|�N+��	�֑���C���8�"~h��1�D[�3v��7��R�0Oj'��6�2������
�1��u9z�'�W������\��B_/9`b�6Y(�@��ך�����&<�Y��T�qA��������Q�xVCxq(ѐ�׉��C�Q�����RCrQ�?[��nY!���HD��`��X��t�6��dy�Dh�"�,�;�ņ�L(H8�{�s�FK��B�2�v�8��&��B��6Wx��+
HzFa@N!�����{��5��6��5��w��A�}ʄf���؟
>Y��5�_��'����iY7�����8��D�֋*���%���*c��O�$���$�م'���e�� ����{[�@��	���k���cL�/:��XyT��%z�p��!�J#��ǲ2���J��Z5D�Ab:�� -� v�%�E~*<�"��zQ�?=��3�̀a^�[3�6��m���;Sl�n0'		V>��Wj�kg<�%Xz�j���SU�_=�6思�X�#����	���)�}��a��6¿��������.�_�Qkps�x�_%�?�������
�S������s������^�w!%��J��8��:�0��L1�\�NB�rԍ� Ѭ��su�s�Y��2����UZ�01���%��Q#�ͷ�S���ù}7?M����5���yZ9�%9c�aJd$N�3rB�B���ޓ������B�����w��Cv{�[e5Ѭ���pi�e�^F���AMZ�/"���~Q��<KT^�-pj�?�}#D�rS�o�e&�rI������}�Hk]~��t�z�;�����^��}�u�ֳ��y��j��đi�?�@�k�)��o���N�[����]�'g�M2�Z�Mj��xiS	s�+N���ޟ��O���֊�����)�|3y��ih���<�wޜ%o�aċaĄ!.!���2����*���Ȇ�H��@Aψ���ȋ�Jf���n:��=zOxc^����`��Mj]j�{f]��Ë�Ç��*��1Z(c
���$3�Ĩ���?h�i�|h���ܓ��}�������<ȥ��0��«;U?��/&"lyqK��h\��|aж�p���%�([*�,l�����A�QM���j�q�d����bfz _�C���PW�F�%
~��ljzӖ�l�*S{=6���^w���"7���Tɪ�s�G���'�jʁu�E�'��3ǣ?~N�tPv	���c��U%��O#�Ѷ�&��qA�k�GZYF��{<��x-&s�	D�O��Zx�	֨�y�%_��S.T�Ut��%��/��`rj�D���=
XolN��I��v(�鞅fk�R�z\�+�7d�E@7>]yo��o\s�]�{yd����u�D�����m��$rx`��<�4���l>����`�Rex��j�=����ſ���a�>2aR�<zf%����n�J�����@�g�g�%��M��6W;�F�!W���E���0��c\N�ˑ^�g�=YE
��h�u]6G}R�A��V`b����������X���������Ա��H��#�F�v�x�>�E�/���j����ʭ	�BOV��9{�,C��4�����z�\t�|U"ܦ��U\�D�x��U�*(�-d�>$�w�1g��tv�p�Z)�%�#�P��lE9������*7%��5boQ~���c{�eڨ�<�8rH�UIV����6n��Q��L2���Z�$������A)���0�� v��4)lC�vy^�ϦĈp��0�A`�UV�H��/�A5|�*�\�JuU<H�� �:_K���&`��cu��G�D1�ݿ����� �������0�i5�ޤޝ²�5���+���ȫ�i16��t4�7Tf?if��j��qq���=�4��@���-T� ��BU����J(i�(ђ�-T��*�Ӥ�v�ҁ�������9#�#���PD���n�9�_���h��G��^��.+w僂C�D�x}@���������5�N@��Sn�wƮb���l6��ǉ�u�։^�y?ԙ2�z�?BX^w�^�_�c��=���}-"��D���?�R�f��{�q�j��H��0>�B���,�s�D�C~���O�<���*8,|���Q�4v:S[u<4(��E�=��GC"��k�RbCo�A��N�#N���ȁ]�GC��z��|g�Y��� ����Q�6B�`��hi$:��R��8�VTw�/�J����#�/&�:�3�ԶoC���ד6褁7jcsNVz�y����2�vK`�}&�E^�)+������� ��CY(R��T�@\RzX�4��� ����dE��Cq/s��:��i��n>��0v��]�Y8�z7w^#�h5KL��C�%vG`�Y�JP�#BJz�|ʅ�QA�E�z]��80��w�Aw��~e`��2�6@�5��`z��K]������V�f�t�5�p$6��TV�W�r3	�@u�L�tE}�,B,��_r-
B�|>L@I��8����F~-%
|_���5q����x�8MK9��/�h�"Mv�	��k�cĤ.G�bG5���j�8),��F��͸.	�v��"����v���������%��0 7����~���Od�f�V}�,�uF�G���q��������dr�隱�K��R<�Ic�W<�n�~*��P�����ɡ~�sj����\"��Wfd��@�ށ�9�n3��N�U��1���5}���כ.I�@�˿E�:H���߈����_�������}������r���)]��H/�N�6ʯ�r�R#NMk�w����o�ڴ�=9pTu����y��(r�y�sz�âI�8����ZϹh����ߔQ���^�%��=Z�	K�&���]b�?���
��Nn�Gx�c;њJ�E [ݱ�U ]x��	����"ֵ�G�x��Ă*�"yf.ni��)Mh|<��fH��%�N�brαr" ��o�+�^�V,p������\3ԃG�y��[�]$E}��PW͟��8N`�2�Eۦ|0�L�6HM���hM�Jm��\ܭ~7�q����WU�'U;L�/9��j��������Ya�Ϊ%��;��rbd��&,1c����%g(˞�Y=��]���bT�Z�Do�,o`�$��Ɏ�2Κ�G�Ҵ��*H�$����I%J�b RjVKĵ�ոC`<��I�)�Q)����`(��IP�5�Oȱ�T��>'f�����w'�Ъ���-;�N����e<����k ��O�Qey�za�:�N��,��{�d��8�A_6f��L��|�~���_*cE����8�fWI���L���,bP�?˿�g�����ɂf��<y�dMC��}�_��2�N-�E�qٗ,�.C*3��]F��y*���"��]�7�<  }�!����}�$�w�Ud��Us3�7i0����L��h����c��*����q���eK&A��*]��~xA\��(B�J��}��Y�q���N�$'[':�?��1�+��y�~7x�u���$J���gj�t�z�P���+8�3�vݢ���4��g��Y�
�	��.�%����A')��9�GQ�� ��S���ƃ�1�w�Q+cn-l����3��-z�/���ɔ�N��4��B� e��&�gP5V�H���(0V���׭R�Cc��i�3g�E��i{��
c�q�SF�M��R����[�z�Y)[��sj��͈��ja"��������O�x�͗�����s��%��p��>�aM�y8�]�z]M����h�	�Pj���6[��5[Y�4������9����%-��W�A�����ߐ���Twx�@�� Z�G��kRM��5�' �m�jJ���C�DI���-�*vL&��)
����_��AZ<�&��mǋ���50���a�gUF�a����!����t{�!�u5��ԗ���<�|X�]ʫ5���b�v���(,�ۅ����A�𾜠��A���^�L��X�!}���� K�k��Z>��K�|:��J�p�~��L}VQ����aŉAi�p��3٩ǃ��;4w�S����a���q�G���sUy��j�o3��1(�>�Aa� B�����х�z�OE�z��O��/��fV��y�0(1]U�x��x<f{�>�2�wR�ZV�P�MrK��'�ĥ���qP<lǋ�~�5%b��k�6���EՍ�=o���=�jT֤�+����X�9-PC�\}vg�w���_G]�r��		fz��_�'&P� f���ֵ]}�^7#~>���58թ�O�~';�9����_ �4H=�?g�y5-v������ե��&�ə]7�:��D�M	J��?�����n�C8�Ӥ�_1�pd$��6�C<^����h/��,o�:3WC�Ai⡻[��/�������$���
���H;���Ҏ^�W[�|�}�&z��O��P�
fJ�x�t�wDH�!+&b�k,Pd�I�ly_'��\g�>�|�`�y��Ks2��b�R�r�<�Y3 �2pjBP�i9�L�o�+�1���a �}�*Tx��n1؅+���f]���޲����3yw��e�K�߬ ۘ�ϫ����|���<a��m���0�m{��){�e�V�F9��@��g٢�'b�<n�;yR�oN��h���}�-(�'�����ò_���-���Z�Sm��	���Ԃ�x�/O� 4Ϛ�>
��d;���0��zE��t*��З�I�^w�ܯ�٤���E�<`���+ ��P���K�F�l3���Q���I�ȱ`5�Z���<��Cf�Z��8ׅ������%���,���-^CQ�S�����r��dq��[J�~�����yFW�w�(���8�,��$:�/����#*���WZc
1x~�푨F���d��^7�'�N���Ȏ�������63f�&��Ƶm��):#7��ə�>$�_�4�9>�NfS�䙳������z���yxZ��(��˃@<���#�!��������\�I(�H�?g����9��,=�w�u���K��O��##OEl8#���^����~Ԓ�f~=���U�.�Ҿ3XP��,~w�=~o����N�>?E�����b��Z��pVj���N�/��9wf����b�yu�䭦(��5􎖤�C@tA`&��F��0��hw5�+�Us���а���ͅMlb�9�(��H*��Ӟ�%x6n�̩��Su4:��'�����ΰX[�}�̦��s��Z�_!}�o�.����_ңJ��Y��q{���`wd��@��s��i���h�L(ۘݷ8n����M|T���~�_PZqPc��e��r�_��q.�͕��Y���SՇ���A����:o����@�R}��(9���%ρ����ݡlLŋL59� �ӭ84
PAyh�c��b�@5fDM�=�`���ն�+���]�/[���i�-��Y0\�&���|�i�'ږ:1��-aÐ�����/%ԊՊz�#��hV����ֽn��(O�k��ԗ.��%j�Ga�J�6=P����(��5���<�wl�)s^�/:T(�T`��\TP=�\|��x��pB�/g����r�H�$�ؿ���"���ԯ����e�i�`����	g��{~�o�;�c��vJf0˩�(͕jY:��ro3z�l!ȤO����W���&k�fO��M{�$#WV��.ם� s��$vmaw���FHہ<�[����3z��#nAh88��ɗ��	�D���>l�}>rO���q�3�O7<�ų�ykό���D����`�-�'e�0�6�A1DltͿ�����={?��I?w�Es��T��pC��	��|r9�(�'vX+t����DIJ�D��I��W��[NP\C�%Fj:�}�̩(�)3hO	J�b�@�ǿr�H��j��H�*Z�	 ;�c�n)b`���M�8�n祉�c��`{��ֽF���oJ}�}V��B��P��u��\w*r�;�`���1q�"��m��g���s݈H�qt�]Nz̗XϬc�2����R�P/�3�{K��j?��}���OE@�d��
��O�7ܜ�6����Wg�k��]q�������nA]�3i=-�_���&T3h�bM�)f	
����N�>�D~�5���/
s˝�qK!�����q#r�N�x��Q�X��ގ\�������G�	������)!�4e�n�GƖv�gE�}�.e�&*�p�,Q}��mGX���{'n'��p��4�7����wPg��P�>a�&BrIDH{)�@���ZB�",�S@��ǳ�J4���&�|m&Ǽc�
��4δ9P��N��r����ڶ�Lf���L�+T���ȴ��N�I��A"�]�_��E��u�ξ/7T�a㝙������L�F9.��*��
�jWxZT$Xf.��;0
v�Q�<����k�j�H�a�!��o�]!bY^3~�Hl��LD��_1鍭��k<5]�|)��orwG�9?��Z�^F�ly-,��M;nv:�C�k>�9��k�#�'��70ShޱD�`�RNU.�`^b�|�����=�'���]=��l�,Ѕ����!�2&LK���+j�V�1�Q��1������i]	����р6km!�K��[X,������{���엸�k2�ϒ��uyE�ɗ��n�:�����#0O���������t����܇T�����_�ԫ��1��&SVtqL�^��1"1��PH�n��D]�S�%�*t�DZ�3�"�zv��Կ����yur���ަD�JV��#��C�?_g&�i�|�2jjF���1t�������1���g����,��mi��#g����S"uB��[��2[�$��,��+���|�S4�l`mp�"�`nE���'7g�qyW���+"/ ��Z��2����̗ؔL�m������9wc,��0�&��aT��8.6��D��F�i/�c0�n�#UB�,���dV�����ܠ�sy�?�����]|��/�57iߴ��^����5p�k�,��|`j�07�Mfhّ�~^��%�=�)ٴ ������8!i����ZfSS?V���1�wE:�$*F�qҥ��j��|�U��Qi��ޛZ���h�c�/�!���G�p�ZH��v$�fYJ�:Ӿ;
o�ZR �������mb'��Y�IB�e�G}�R[�鄋�hv�W�f�8������Kź���L�&�s 7v"�A˅c�,��	=$G}�	�����ش���|�1�P�(�ײ0�ڕ��I?M5�w�>O\�|@<�OPR6�
���W�G(�-�Jl��VJ�f?�Zj���Ih�ӭ��
�*kv�cp.���%4���H��|`�"ؔ~�r���xGZ��h�m	�$���5F(�3������DdբQrQC�������7F��D*�dh��s[�������{��˾�1�,��9���=�l��>�����߯��S�����^��S'��tG�&��9�ŕ�I�uWGNhʹ�,��:�{+mx���|�	}�y�/��Q���h9#ߖG��sP������a�.�V 1�bkzgip�W�Y��3�g��UbT�Dy5��@�&�"��/�l��	ǖ�f�������U�Q���1�ZoR�3:�iW�к�<�-��!e�J";D��m6E�n�EE� ��C
����oX�<�� �%$��!���5�'O����G[�7���,;ƢM��ǭ{�u��nZVm��>�K��ت'��Ju�j�������d��ܲ���"E���/b�����6>�y��\M���u���$o� ��d�x��'>	oӿx��8A�7²���Fbdd�h3iY�Yd�����L�$����Sx��βV( go+��~l �����[]�g�-���<LqK(_��!	����%�It�I7�c?)�r>�Di`�K���b_�j��uj�����M�j�k�#3�����,c�=�m9��g<�ĉn�+�j�!9��Y���n��w(�bLrM�!q����T͔x��d��`٣B7?�$��@�.҄f��,-j��x���mq�����5V�' K��|;[��@c�k8���6��O��ɓ��~���"�g��������]�N��-�؈^�w	{vϲ�D�2�1�ܙ�/N�]�/�iRզ�����P$x�=�*q��	h���x/A�y߈��$�^OY#l9yd�uX@�R��6���	������.#]$V��,~zǵ䊣1M�V�-��� �eI%R�ZK�������c���m`��i��ձ�I@<bcb����l%�x��@��,+Z2	�,�蔇�Ŀbd+�� ��y�ӵ�R���E��q����R������6����O��f���e��co'9��( �C%t{\Z�!-�D��m�7U�Ra�ũ�ʣ���6��:J�M�'ߑ6m�
���^>+=��Պ௖t\Z�=Q>�O��([R��G�����cɼ��ݫ�I8��K���
�z*W��(�M�
�~�~60a�B��c�?G��8އ�'Nˏ�ix���U`��A�H�'�e{79�1+�.����ki�A���T� ��s+�rT�6:ȁX>�@�/�P˔���SZ�cՖF�����Ͻj��L�8��h���=2D�L�o;�^lP�A`8����Թ�#U���!gN�1�Y,�
�G7L�Oe7�W����S�+�\_����2��r�H�0��i��/�g��v
��y&;�G"T^~�0���)u�y�=s�>����_Q�^�z5�~ޝ��?��h�Yz�����Z�s��$9�Y�a2i���ރ�ݽGpj�/\�����bY���-͏��֑�����f ���HA�\����X�6:9Jw?3;����h����7JH?,/�a���̯���5����a�P���|ZFϷ0�(N1���TXK�(��D�I�R���/�[���M�.5Iѕɉ�,�P1�̛�(I[��.1���ϩ�'[�N%��Y��: ������4ŋI���Z�W๿_g�l�*�ˋ�޼��2��� ��d�a�]����=������ �Ю��-�k�p�P���{<}~d��a�7�ոf~��4�RS�nװ��h���4	Z�J�7q )gğ�N˦OX���,.��p~�/��;Lj��`�|���&�u� �����X���#��ܜl�f��w�{�~-�9?�ֻOjMx<}6֪���;��b����r��ȍ���Ԙ��d�;�&}β��Q^�C���8_bO�Lu���d؂�&0Ӂ�Ӫ�F��zr��K��hdt�dh}	u���Z��s6+�i�Q��.����U�e�lzMc�F�@i;��s�S�/��h��e3������z	��A�����c�̸F�&�����j�du����E�:��HZ��b��̈�������{yo	�|�~�����`����?d^�����^�{_}�N�NhS��l��gĝ�\�t�@y�W�j�;3��v�祣�<�5�u��z����F�꽋�I[��Ȭ��p��2G�쵋��<HS_�Ȕ�+l�XnG��FR���L�����-[%[y`HE��ȈUy~WN�=������l� ��Ȇx& �z�,T)�%:7����U����=����@Z���UR�lz�%9�	�4v ���|9̬����몾��bi�e�gBi�g��Ĩ�8�����:Ǥǉ��0�F���Ñ߭��{�$5&�e��~Wd�h�8U�7�@o��3N�oՖN�4>���4����f~6�Lw��N� �N$�����n7�d]hTt��lS�
��@�݈n\��Y�DX���_���Ρj��8��O�n����������u���qV��8��t���Y�R�R��ޢВ\|�VԈ�`�'i����R˦n�Y�Ȓ�,�x��q��*�O�Fb�aT�5�bV�D�q��Ԕ�w�Q�$��Qr֥�v/hR�%����W� �>

K�d��Ћ��PX��$� �
��I�ģJ�O��km1��C5e�uD,Z�dX�0K	;�Z�F{���LD��UB1f�(��Ŝ�6��d���V�L��DP�������k�TER�tj�5�0�ȿ��N�vO���������*��3�����}5��Ed{���ޯEp����
�%�պ��5OWNmE��7���j%��M�Ơ�y�J9W����#{ݟ��B
(hkO����h!g��ur��ö���_�}�o[uE٬���	�y~Gm�X,e�)�RG�-h�54����q��AUZwG��F���[1}S��Z�p	�Ħ�Z�����<s�Ӿ+=�L)+�o�1�M�[���G�7jx�)��bWT�T@f��I�^,���41��:������ə��ս�F�Ƀ߀�n�ԏt��D���k�,��u|�>��=ߛ����~dAq�]�
rmI���V��%�I����vl�Y?��<�f�ƈDh��I��6�]c��p�㿾���.��Z7A���h�ж#fŒ��6��Mp=���t��őm�Q/�M�����!��Y�8�zR5Csc�H<�aK�F�%�.n�{D-L^7�w�襇	����1�H[�-ׁ�2h��l��< Դgj�4hͨ�6��.o��݊6��`鏒���ԪBl�"����br�a��ʢ��@��b*!�Hx�?��*3��D�8H4���t�|�XRU�!uy�2/�a��H�!�Ba
�V�+���n�hJ�B�C�h�a��i��٨�e�G���N95�4�����ϣ���*��j�����I�-l�o��m7,�v,�����7)�`���/"�Y��[h_�UїV����>+3�W�����̩k�����5A�~���i1N�^�����9��F��w(��A�4�TO��f@�ef���*�������Ou�%e|f ����h>Ǿ�#4N0�"�D)�n[��O]>�H2��Ys���:s�"��ƙŒ*�{�`�kL�e�J)(9�"�����p�$�(�M���Z6m���C�a�#���*�QH��(�p�A��bT|�C��{>K�����0���3u��N��4UD+�~\��N�p�d9�Cc-���-(�7�q!�p��|�a��ݵ+�΅�d_)��ʧ� �iȲ������Js\I^�S�JS|��V�b��l3�㢖�f�!\R��z��
��ʫb�����q��OTB}��b{?���_��&��A1v�!���a^?��n�G���Oo�g�
�+�K"d���cM.�̶���8�4�$���pMJ8o	�c������~6`}��/��/�!�mi`��u'�F
�m���)�yT��`�:���6T-�����|E�+���}"0�Z�KԿ��zL��=�#.�q��ۃ*Ԍ�WI�s@�d���l5V��wOY4X'�Iz��Dr=�� 7�R��x��=;6�� V�3/�#!P�N�����<�-�E��} ���_n��?��~K��_���C�����饾o�������2�D_}�ϻ����7���ƿf�e���e�z9/*��B��@���Xm֘w�::VL�Fm1��.q"��}@�G�ޡ�{aΞ�:G=�q4�₸��F�Zl�Io��{�,&[�PB��_��r���v=XC#W�:�>o�XO9��?W|֝��o�?�f������+)a���tM�M�&褙%VZʞ���4ĊB]��0C՘�Y3J��	�/l-;����?^s�!��'۱� E��k��	5��P�/��
��Y���_�L	�߮���7���_�65E� ATvM⡗�/��'0�Z`��3�9��y��ǁ��,�,�IJt�#2�q��V���pWlҨ'�U��EO%���B��i*�V����m�6��s�u�x�:�S��\��*�=��[��sղ1���o�}paS�L���Ĵ .=|��5��M7�إH���3�'������6�O�Q<=";>f�h��c�=�G��-DQLϰaZ=�͍������̌�ghjȰ{�q�xn��ð$��q�􆺪���e��J⡙������P��vu8�l�g��Z��4ۉ������2��U��3��T$�<��J��E��8�^{��F�w>3&�2����I--#�B!=[��Y���Q���B�㓉%/�꾟�+���ì��u���ϓ�l�x�	X�7���x����z�mm��>���&����@e�҂6�t c�%��ӢA��,�rJ)>����b;ߓ����Z@le�����X��h�AE��3@�J��:>*z��͕8��Ckm]d�H����*�?��]���4��r���B[x���N@������lX�,���8���Dv7��!�Јx8�jRj�!��_
ݒ\i_�'���$��Е�V69U�`j���ϩ���!]@����Z�׏�6ժA���zsX55�أ��'��Y�	֮���8ƚ]���AkbMt#M�)��m&�W��V���Ɔ9�kG���K��2=��#�c�`�����E$+�s�@����61���u����S�?�X���|����{�T7V��%r����O����s-D�+��C��r�7Ϥ�s&al���	$@O���V�fR�)��r�����1Q��07HFL*v��$�i�8T���S̒N�*Z�XlznD��)�P��Qk����B�H��A'Y6�6�X���H44�4�%����X��X�G��"[��t-R���=Җ�h��e��nGB++�h����1�wʧX0;��Y��|���2/����b'c�#�Z�l��̘3�L�4�{�r�uwp�CϠ�;��4�!����|����}3>O��cj���bh��7e����n�͟^�2Y2v��ܟ]6�ϥ6^f�e,\���o����e���\H:��p2���j�ٵ��W���(��E�I�|�hI(�D!���鈻d�
�<�N�t�)X@������?�D�)�L�[$K�P���b�F&�ӎ/�=$�k�ߦ�JFE�g$�$�|q�d3�\����� ë�Es7���Ibl�����R�l��-��텑�jlA�J�u����4q8�z��q�hD���L߯�ٞǶC�V�fC6Xal"ٴ�%lʺ],e�hkC���j�+u��#��ɻ�
�$�q,-�:�� 8�6i�̫���n%����*�ƛ*J_�D���
�0�]7	h3ęS!�����`�����򌎍�z���KB�P�R����1g�,z{f��+V�噥/*VĴ2��R����NE�AFO��Z���kA"���*T1��i-���A�
0���\:�i+Y��-Җ��t����s��4�YKj�i��1iz��!�6"��5F�BF�m<7E�ҕ��u�X�$d7��4z3������֨65̌�olPg�Ey��^N@#h`gs�+.�n��$[���[��P}c-�l=�o��	�F_cޢ���e�n#�P�t�J��^z���N��a��m�ȣϽʥ���f��w�����O���)@�|�N����S�f��xSV�G7�s������2�<�7��'~�y}9zK�ԫU^}�U�f�`��5,_����h�"����o�ݢ�����_I�0�ZS*�Me�NIv� �@����P�*Xm3˦��dR@䆴�����ޠ$S$��7J��A�m6����YR��X�r��:i����XO6t����eD�NF�<�
k��<	��p%��*��ݑ��P�A@���I���RmEG�X$���IƉ�͐���:w"�2v"K6l�����`��b�u��&�1���.NZ�Z��6=ż8VF���K�kI��z�(��nh��8GX���M9pq���+"���a\��&�y�h?�Q��NS'�˩��M]�o��j2&��䈸V�Q��VSe�T��j�#�U(����d҉�=%����<�{I؏�%"rM�5F���x�b��F]AʧN�:�#c*iy��"��N�3�m����bZ����f+t�:i4�g7���գFy����Xv���W�c!C��14S�0q+��*���t�M�)c$�!�"R��|�^+X�!qǢ��T��Wk`xM2�IKk�M=ebx.�p?�gg���x���Y��������8�z�~�6l�����0w�<5Z��:�����W�@�7_+[dxx��?��N8x��ޔ��7�Z��e� ��m��~}��~w������ze5����l���ٝ9�׳�7�y�����
�)�|����δi��Q�������~J�g6V�@
3���d��:��)|���jC���ne�v��֯y���ة	�S�/�i�6�x�- *�J�����ha��5�lXM�ZQM�3�m��ic�!O�i�H'�y4�^f��ȥ�y��dd��9kg�tw��'�&Wt꿣$1x"�-q�����CP��T#)ѧ���(i�F�V�K�� 1]�*T��G��Fa"$80�ܓf������Ԍ��O�3��
0jI؛c&Y���/rl�A�T@M��s�iJ���#ꄭ����Z47�DΊ8r�	I�j�D�HN4)r���J)w��#����e�)뼜�a��ol]7�`�k�`�Z��U&*`I�&�4�2塕��.��brNL[WN��0S�̻��I-�j��QQ���hy�Z+�eRk��H24ju�f٢C�����H]��,�h
#eh�f	�MFOMw��{���DaC1�A�$�T*W�����4�tIg3�3&�� �7^�K�ܗ�:���NO�t���jMY��:{Q��b[3g�!�M4�`�p�3�>��Q#׃�mcdd�#>���?t��o��ԛL������S+p�o������XJ�\�'ܑ�}l7�2�g�q�}���t�V#Oس��Ma��9��O��Rv�O�4��-�>c冇cfU��&@)K���b�L��h��|5����ky��!�h�u=�9���*X��oҹ.�sRP�>�V���(��U|���CF#�W�@=r����3n0w�^_�B�3B=ˢ����g-�%P !+w��3
��I��f2B�hm�F�'���Ϊ�� l�Έ�&ɾ��E��D͊q��Mq?!beS�4d�t9(]R�����;����3'Y+�/�3�F��l�qL��R�%�`i�v�dL���Xz�@�S"���}S11j�&v�	���I"�b��� 7���F�'�>�l�#�I�uJ��l6��]�����ک�H:��w�@A��K���$�X��R4;N���5H0���0��o[�T���:ʵ1ꮯ��
C��J��:wC�_-_��\�Ӣ�I3:>�f�8Y���~�:��(��c`PG���ww�md:g2�r��ǈ|���E�LXL�mr���Ԛ5JE�&�1b�FU.)����l����t��93bt�k���쵤�i�Kv��vx��X��B�}�y`�x��l��Nd�j-X7T�;߻���&Va:F����?�ك�9��[˼o�5����bh�#���{�����G"�`lh5�z���(��dm���9<�ؿ����������EOW�aH����|���q>3�e��*��@	�Xw2�cr�0���ƒt�S(InU�9Q�U�=D�ZO�
�=ó���I���I����I����R��J�V���j�\���
z��Ի��Z�B�&M����?/�E���Y�r��
L�:�bμ�d\&���J�M
	U��D��҂(7Mb��p6Ki?��Roհ%�w"�_6yq%	@T O~N��L2&Rap�<��&ECiL�Uq[~b{�e1���d­I���"
\2&4*FG��j��&�V�T1��$g�c�V��b��k�O��E�j�j�ާ��O��L&ʨKuO�[(����ؖŹ���i�D�Ng+��͚,RR�K� ������dC�n� H���Z����|j�^>���lX�2�:�t�gy�'�5s��Y�i���$3���q&��q���3)����X�s����j���Z!�������eø��=�����X��Z0�RǑ�n�d�y<��r�I�S�d�����F{>����ا�r��"e��#����3���g~�6��)5�4c�en��V��5g��/[�"�v�	d��,���_��t�\H`0sEh���)@���dk���yk]�w��\��G���_��#6ล���݁�q���:EE��8��4�*�.R��N�|��~ҙ4�6���ȫ���N����^�%�l�"��$����G#�$]� �q���>F����b��20I��V��#=��cl��ؓjeTm����,C��*�T�s�؇�h'�l��TX��#�Zk�S�%Λf֤�Jagg���Ӕ��tF����|"W�lg�@� �HB��e�t�FD{[�j}�#:����2�t)t�I~N\7a�&�G�Q��W�k��:�aebr��j�R�ߓ
�>�&%������|�CI��*q9r�n�R6�d�&�X�%�œRCM�M$.(C2Z|��6{��v���S�0�&�T�ЈhZ`IM� ����0�b���a�a$쎌�6V��\'y?	K#z���0C"��`N��+02�~�=p'�8`>�<xfu��#Zn�01��y�b�"��,�\�+V���I=	KJ�a�!�k6w�|^x�%���
عV�i��з=g\�+�Ӷg̕��461yäY����вixUr9�b>��K�Ȧآ��o�D��~�~�b���1��1� MtZ���Y�*G��|�#�)��d�����2���{`�~���c�ڐ��/�V�1Ll0��<ccc|�mu�G�}��!6ubo��4o�K��8@ah~z���ںI;c�_%危�N��}�RV'
�*�W��"�~������G�꧿��L���EL�I��D���$��F�d��+-�p�P����2��מ!��8!�ڰ$�_6�&�lLCB�̉����1���g��/��<��>�N��E�}L��o�����|�qz�#Rn�f-T,��`E���.
]���QG�?:�k�]�%���z�Ğp,�۩��I�v�0۞-ҿn���q���]|`�=��]��t��
Ө7��:�0T��'cM��tt�{�=y~��,Y�=7�x#�B���a*0��,52���@X-R��a���D{�1c��y�U�-~P#zdRVJ�LR��gxԼ
z�����Gc���a������ˊ	�V�;��RQ�CR G�W�\4�C�(7�t�r��{/�Z�|��������Qaw�JOx,�j1=�+�i1O=��Fe�����~�������Y�R��l���F��0+��J�����=��{�g��+hk렯��F���}|����(�e������2iUR:o�]��ïs�/���]<���洓��^`��Y�~��4��`��u�x��3���{�lEet�����b���j������ʼ�>"S�Ao['�V���*�/~���ݝy:�r
��y}-��^����^��~;�=���k���h�YH,Iݎ��ͪs���my���_yg|bM���q� ������_>�Ǎ����f�{�'oP�٨�ّ����̾ϝ+���z�~�x�Y�ǅV��n;B�R&�$�L�&&�i�t%}�J$*̈j�Ak*���IAc�ru�� Q�$�D�� R��hC�eLҖIKJ)͘Zm�i��̝9��Ct�X�H� S�O˗�G�c�����X������5QN3M9r(��d�>�p�!^l�-��=�6����l����'e��uM14"�6�=��΋Y��r��f[��e֯��XE�`"?Eq����K�t�6�Wh�(���;�����q����[U��!�Bx�"dN���}@#Q��Z���A}��I�%���Ct��%���Q%��l���bhRbЉZ�^������m������v�z����6��T��$�� q.�I*�\�tFg��w�{�e�]w��?��K����#�P<\���R`�or����V�2Z%����;���p���H��߄�5��`������$sexo��Ɓ�̣Z�)�F��
FFG1-�lZj-4FF��Y���2�d�����ѓt�Eq��{Ȥ�_���y;q��+���֒n_��������t��0P\��ŝ:Gf_^������I���� ��*x�wi��=<S��>��P5j����veִ�u���������̙���_YF���ko�w?�4v���o�+JFT��M3>>�_8dJC�6�l~'��y']ͷ������w�u��3��C�zX����uSj�n����!�<9F���i�1�b���bl2�V�'���aio�C=��q�
MӒ���F��l`�����&YK't�n���z��t�K�Hi0b��2�.~�&5х�b6���5��J@�}�աD���bj>��k^_����"b�F1��*;ǚ�O���L�;=���'Ar"�M��&y'O�RWVn�1%���%��$:�-euB��eD$�q��x�q�8j<�d	J����ȖDkҢ�j��H*�Tzp�����8eIΏ0$�k��W#SȪ���)]z�Z��N��x�Tb�n�e2i�&�	��k���	p�d����<N��.����N�U�/3=k2���L�	 � ���@ E@A�X|DEY\^DY�l!� �@B��L2����齻�:�y��]3��#Ͽ����>U�9}��\�k��� ��F�t��K�/�젞 Z���	�������e�s~�T���IH���]'�'Clց
�k{!�b���#��;_Ǖ�|����U��Z�&��lQ��t��lߦ�)�@�x,����n�)��#��|� �JEM꯴R�*�vlk
xU�e�V�@B&��9��Ⱦ~�����̷��C����!H�_�Ds�4�{�e��V��Xdbb3�O��Ƴ��3�]��Zar�4�x�ly�{�_��9Jy�"�gЦY_b�����FL���P.f�x+kMn��>>��`�%R�V����� �W��y���/]�����>��[� 4�����&����}��?��*��&鰩�����7���jc���+K�9ݱ0%V��|�\�@�� ��ݞ�ȑ�s9)O�N��Ԕ�ն��MP �4��MD��8A,�!�!%��1@��rEU�+ �3P *Il����_M/���6t	YK�^+�����+����X�'��dt��+��.z��\�0�jU�P$�FBؒԁ���l����K	�h����.�[�	b%�Xz�^ �*/�%���iq"���8fM���z��Ej���=M�0N��r���i�nF���c�L�!H}e�`���(��l�:YZ�3~�&p��,C
5-����4ѝ�z�~Y�����2ԱE�"�W�)�D�j�Y�ύ�z��W���L�}9?fR�(��:_'p��2a3�w��X6Q`P[��Y�n�7_�4f�®��S'_)q�̤b���=c9̜9��@E�*q���֨V�4����j��
;�����Yo�k��\��Wf�]S�j0?���S�̜�rL�Z�;���d��o��."��d�r��\qͅG����ȖA��p���j�k�������y�;�M����x���Ǹx�^��߾�W��Qf�[Q�̡�"�<�������z�8�hu<V�;I;;��)��U�a�ߔ���8J�|�˞��m/����[��������I�i|䏈���_���?���sI�t+T}�TP./�P,���s����sj�R6f%��kl�ihq����R	a�	Y�X�	6]�鍦�2�z|"�����lV)��d�X5�����B6G���Z��|�ʪ��Z�M�:N�c�i\��.%�
yKt�N��k�غ���{�φ�a�6�P5@�Ȩ.�X���u;
�$H�k�&i�IU�B�X*x���E�    IDATzN%+˗ 4A�2J#"qn6�0d��# �u�t"�al��(�d��+L��"����#��(��� ��$�:���Q!o�Ro��QΙi����^'c�·��95��WY���J����G�]��_�	`�t.X���ci��{�Gz�z̉;z���~.W�R�z�O~�$���C��)����L��fl�b��H�M��Y^]f�舺^�9B�\V���d�%�!����Ţ���뢝�U�_7�/Q*��;:I�Ǌ�N!�U*��ڔv\�{��+��'0�1���R�xuFu�����c[Љm�z�w����������9gg�)�\Μ:J�����5>��/1�V$S�P̟\ۖf�m��Ӏ8jDM�y_ ����1ݚ�-v�6������( �+/{�����ݏ�4�/��X�ಱ+p!V���t�S?��_�~ahϏ߆Lp�)]5(�CJ �`y�-Lå��)J��Ql���E�׋����\Ѣ����R��ר'��l��і�d��w�j��T�D��z���-�@5iC��MJy��k�����W��dB<�&|�K���)�4aT�.}9>���$GG�B2="��M0u��SP�4�H$�8��ޞ�V@���N�8!��)���'�izu�7e�@3ӣ���9!�d��.*�vH-K��TUT��� ',����I��%�ͤ%�F�L��@�|�D��MY뻭:�#|K,ɨ!L5|ɹI2h���I�_��yD�'�!,�@�OUE���T%H�����3*�s.���a��z���%M�j��o��P���1��9�7�����H��8V�Fc�%��#�T(�~f���*�[�<�����u)5ٺ}�҈<p��+�T���+j�7uz�15V2X�_�P(���YY\"_*�n��ho��1�Y����yk��=�4�^	�`t`��a��d,�����|��%>�o��P��u��}�k�yǯ�v�~��8����Kv�c�޽�t�˩��U�^܉Un�Q������̶G����~+]#�?U@�]ðt�(U�'�uZ͎zo���/y�-S14�nz��nhh.��t���� 4�Yah��_�;�?H�%v�U
e/�c�a����Z�rbd��U t�mb��&SIJ�H�{L�9݅4�j�si��*�BG�BJ=��u��e2�Nz�U��	���Z��R4���n�aa����$��iU�������;&[���J�����cxt�N��HC)G4q�E�}C`\���E��~E@����K1�4�~30�u�ɱ�6�S�h��Ű�B�1� W4D�f�.����l��%���F�M�ZE�(���W�'	��9� ��M����iF�bd,"����K��D��F&�+�E���Q(���"q��������Q�V���q��I�"b��(퍖 i��nG���[�Bh�R4�X9K�� �ޭꉴg���\��ym��l�]ʮ�ccD�t6zo�(?[y��Z���G���)��N0u�v�FFT�B�-+;VgO�26:ʙ�)�FG���nc�9V�묮4XY\WY6۷�R���zc��8�J��M��`m�:��3,b��YG���a�k��w�ﻃ�6�S(��}�k��x��w12`��z?��z�]y)[�6��W��_��ZW�\����L�|������?�#�n�I4t�'K�����}�|(}O�bg�9�T��Y��rp�~wT�����闞��-/�ֻ 7ԍ���� 4�Y��Χ������� �.9-G�J�Y����)������2eMR��e�Li4[$���d��q����I6*� ��)�TN����j�λ:Q�Ή��{\C��	ݮFqh/[v\N��Q�0�r��wi��f��!�KoP��&$f��Mב-n����]WbQ�	ɘ:F\����"nװR'��)�����_���f) ,8�y��<��Fi@Y����p��������Gp����n�%�ce���+�j,�����hv�P�8�K"=Q���kt��L�/h3�iՑ-$z�0�
)��)8)��YN}M��dm�^z�:1c[�Q��N��qSf&�^=)e�F#;)oǋS��ũ�)g\F�9z��JCC b%T��,JES#4^/A����c����5*(�?�޾^O�cyΥ+�1z�^e��k)Y3�\;�[^�4�<��ΫM\�Oe���A:~�VcS�l^�u���1}�|��>��Dp-����6����^-��������K�R�/S)�5^ik�*�^'R!_Q����&'�y=_���w�����y�#����3P�����+�����%�<�Y/�o�����x�����:�_����s�;ma'�D3�u[(�i��D���F�%�39Š�p�Plj�ꑒ���S�� �+_��}o٨>� �Ӎ���� 4W�Y�}�����n�vnh�z;�h��eƣCm�,7���-T����ة)W=�� ��A,㤞GF�,T%N�ǹ��F?h�䬔��s�G�Z92F�Z#�3ǹh�u�{%�}܌��Yf��dui��:���\+��'��;��V!r�(�y*Q�+gh����X��;�5�0�؎k���I4�)��=@fɸ)]ѹ�ٰ�-Ku���6〙vi-M3?���1c׊-9�9���H�N��
�ot'աd�#t��4
U����i�rlD��f(ncx�.R�D,:���L�/�fu�83B�=a�TB�N�R�����H������{I�SJ��3��&7��v���39t���e����<A�u��C'�$	~S�F�rz����������UC��<���x2���J�ω�U�C�(@�X�j/��P���"�g��a����R��)7a�.+��[k���&���
����*\y�u��ﾍ�/��J�L�Ϊ�����<KKK<�0�x�+ؼe3�?�8�R^�_��m;}�u��
���2{f�F3"7���})�Sݹ+[FkkĵS���Of��,�f�W���}���K�����M���NkF%�~�A>���`�e�%(%��M1�+mU*Ţ��Jx�7����$�6GƁ���OEl��.�sζ���x�7�)/�u� ��5��[�~�g}���^a���qj������Ϋ^�|���\�u�j1ǣG��V������}���P�E�~��"2U)���+-���x��+ZM��*�l��1{�Q���J��]�2~vaX�i��Y'e��Cx�i�Y$��7t�D�3�
�k��n`�m[�S���5э�����e� I�A	в��,c�ﻘ@sH������T�#���G�Bh�J�����ܕ�B�՘?�8��9�=¨�m�d$[&G��n�*:��{��W�9����2'O<D.�cb��2=��Ц�l�/��Q�U����Y[8N֖q���HwQ�m�+�1U������V���QZ�G�U�M��WCv_�q\����м&*HP4F�lI�R���E3a
��*+d"'�B��)�J�VU�l[#c�P���2�ى0W,�2��d��J���u�tWN�++��ˮc~�a����;L����c[RyP��n����9N�P!�������?}?�J��.e~~��}����|��T}�e\r�.�LO�������=9vSO��Z[�Y����QD�PQLI�ZR�Il`�v�^ɯ���p�\��@�Bc�1����jO��1C�Q�󟿕/|���������5Z�e����ٲs_��I���G)_DC�����cҪ��[\�}+۷l��Su�*A�~����rTQ��U٥m��}��Ϋ��s����\��O�.�q���+����O�.����?������n�sY%�5�&��y�s�獯{%�1�?p[�o&�s���dtd�C�8qz�w��/8vzQ15.~d)1l��6�@���$��JvF����Z{���&��j<���c*�.5�*��D���F@s�1fO�G_Y��l�/m��b�(�ڕ��T��z(�J�ቫ�2J�n{���*�!́i�Ȗ��Y"-FFƕ��p]"�P���Q��I!��y�HQm��-�zq���m$ئ��oZ�u��K�5�&�ģ�:��r��O'5)^���~�M@h��av�a\��X?�1��ӳX�,{.��V��,F��&M&��\@���>�<�Z#Q#���S8�
���iN�2:���S��NbK�_l�?����4:�f��a���v���U�a�X�	����p"���� C
3p���	-�p�ʑ�%��'�/��bAۅA� ���Vd�)ܝ�J��hpt���!~��v��2�z�8\��;�v¶�d�eN<~�-[��`GѰ�V�T�w��>>��/����
_��y��������y��}��~�(��_��N�����Y\��Y�z
��.�L�Ү�@�P��X�Qo,��ݎϦ��e��k�����k0s��iͥc�p������ؽ_�����&���{۶�k�y�z������)<������YL���av���R�y�3��g���������(��>��[�������9�����2���鯼�y����.����lfc��
l ���€� �����o+�uשϟ���+��ƫ�d����G�>;K�\���樓�2�?��j�W�ڛY��[Ǐ]֥��1ql[�P�I�J�]h�����Ato	[���|��&6��<�Nm��fJ����/[,���n��e�F��,�ot�9�2KV�>�-��ed�S)�Ѯ�an� ~g�r�@ڴ�{oDw�T��YF���J�T!�(I�����9ap/W�'��-���`[#)�{�`�K�S����\:M��!�R��FW`�EOB�˸N����O�HV(g3�mcjf�$�0�s/]�B�"�,]�N����$��R���]O��N��,Na��ݔ�:�X�,��}�<���$�d�>�2��r��� C����z��ڣ
���]/��/��'ƥX�o�蜤bB��J�*��R�L�����؆� ��R)Y*�#�J�z~d%�C�W ƶ\쌫���H��*@�/��K���=��`���i�n���m*ohey��/�Vﰰ8G�r�5�s�#3Ć˖�c*P���>���|��� ���y����7�������o�Un��g�뉝�^aj�XZM�W݊ьTe&�|���O�]�S��� �}E��i���=l�wh�N�L'�'f�Y\\Ɖ��>�������1���Ee̼�.�)�">��¶���/.���4WZľ��x���:��­|����#n���E���,������̷���w\���A6V�'���ٸ,.�
���o��t�-��>VW��9V��oy{�W����f������]wQ,����+/g��	v����۾ǻ���h����N��<�e e�rH2)Q�)!�����"@���I�4���q�[��~(l�N>���N�-MS4�x�y'Kl����\q�0�S_����1r���TƯ�-V�>sq�����Pbl�~
�	"=K�$JC�Kz-�J�f�H�et�_�:zoÖ��l�R�yrd��V�JN��q��{����Sk��6�����Ɣ[��~�N��H�1��O����Ԛ�N��m{H�>R���1b���S��I��0�S���(�3� �g�fb���C�w18q1�ӓ�M���izƶ]�Q�K����:Ks��8� ;.ډ��H��pZ	hE�,j	���|�����[@MB��X	�(�f�Nαp��?�:z��;wr��Y\^���J}�N�N�Wɿ�6��q��UOb$����!.?p��Y|�C��G��R�r���dh���3<���S��O��)��>�޽��כ��;���<����=�%���}T%b��>ɛ��=x/�����U1 �2a:�D�C� nR��a�&��}��2��/��|�R��aH��F���Z;�D>�U��b�w�}�;��ӧ4<EKS�j�3�B���':���]�dW����6'��^�"�dqE��P��6�FzA�0�}�W��?�v�Q�28�����-����%?�̟��_��rC�8��
l ��k৵���[���[�Uwm�Wfxë^̓��ɖ��2'NNb;9V��J@�u�aТ�w9p� ku�X���~;���Rޡ�NR�xb���,�6C%n�=u�x}��.����a�c�	���]��!�qX[���֤���Nq��݌��X�w0�[��K.�]벺p��H��dG�atb+'��fm�lVWάBa��{�|Q�X�Y�Pfi��F(R�K���MZ �d��V�ȥRo,�zB���G���&�V������|�V�E'O�S�lgh�"�|?��$	�1�S���ҮO3=uMk��*�ٴ� �;L,ŏQ����Q�p>�#9Ab��bʤ������)�l�k	��	�_r'�p�4YK�<�#;ɍ^�fU��z~�Q��02>F��k�y��(FC	y	�� J���
�(�D�(�$�T� 7��,�e|�0������ηy��^��>�1;�8���P()�.iб�f����m�|�m��9� Ŭ���+��$_�+�*Pt7�>�f�}����߸���_���i�Y��[����^�/���������y�k_�M7����i���/��W���!�HO�Oƕ�e�r���em�N1�#�=:�Ϛo���/��>~+�͚�*;���?��Ԏ�� 7h���E���N����Z�3���p;�u��D�З�h�?�_��k���=��>C�Р�z��#��OƱضy�zm��{/�S�w���5Me��
r}��//�/}��~����O��q܍�`h6�����۟�/7�,I�m��߸��\����֤�&�8x𰲰Jڪ�>>z� ���g>�f'ai�ͧ?�e>��/Qؤ��0%r_Rr�QJ�K�]Jކ��ct���D�A��2���M2�<	�#۰sW�l�4�܉{�R�D�a��S�&�P�vg��Eؚ�U)�Y�6v_z��������Z=`�&6^7�P,@-[�44�YĶ�
�c"z�^�J���q@s~����C�*�T=��HĎ#�N�� 9A֍�����>	�0D'��4	̨De-4�:^{�ɓ�������~�O\��QzU�(�HH��M��'ki�z���?$h�%g�D�u��v24r1gN�j��Z!~�d���3`VI�s�!i�P*2���~�pT,��j2B�W�D���{���kIE*a��{Ec$!}��g�F'�Ͳ���6����27/}G[U6_��1�z�ʲ4�o|�>���J��!rF�����g�=@i:�]_1)#C��Wٻ�
8t���5nx��|�ӟ�o�M>���n��*en��+��]���F)��6>�����/}�j�%
��
q�����͵��b������w��gY�`Z���6O��z*�9Z�e�(��;�G�o��Z����n:�^�[T���8Q1����u�Ǐ����<��l:��G%ZK�����Z�r��W]�����r�m�����4}�c����'�y���/x֛_xٷ.�e� +���l\?��п~���|���x��^�5�/A������Jm��y�0��>r�$J��I��4E������0��1t'G��� OĬz/�ߌ��2�8�#�3!�����Bi̖�]��ؘ�&v F�8�Y��Ͽ�����g�,o��c8��q�R�dn򛄭)�$P#��k)��|�>��"��Ǒa�ZHM��IW˱���S�f�War"�+T�1�54����sŋҥ��;�ͨл��4���G���6����Ko�����f�flqSi$��+>q���c�P��T�@���y��Θ4��X�\���Y��N��h�����oS�)�I�N9�qƷ������,>J>!�������hy�vX�:��>��.~�^!t����R�{���	���9���!h�2,��=�!�g�Α�!��Fh��IoXG�PVWWU�m�TVB[���6������.��}U���h�aamE��r�r�N�Q,UY��*�J*��E����?��������վA�<v���)��)�J�_��7�̎��\y�~�G�F��x�j$V��F�	1Z]$���%�y7�K���߿L l    IDAT���N,��@^�bx<|�K!��2���D	�c~������o�^�s�4�!�l-��p�^^�����U�n��6TEF�y������+�����m"J|6oߊ�$<|��~�?�kE�c��A����%�}�[~��7Z����n��C�q\���O������;:�O!k���y-��Km���>N�|����w�m7�+���صk�/ޏ�,�t��g��}�SL켄��:�D[�VQ��j�7B�vX9s�=��։��a��s"R��Hm���}hN��[7{K��%�fN1<��VX"L�� }e�ř��X=JF���b�cxd���#������[z�I)b#�D�eh�6�.��>ݔT�"�^֊��g�>gA>gQV�2��՘)���7Ly���1�Z�NdA�S����}
Xd�U�b�O5�J���I��iӨs��=X޼�L�
[w\M�@�K��M�HC�&�$�xi�����:'���N�,�}2�%�H��G��J�zLfp+�-�Ӊ]���[��[zH5���+Ғ`���Kn��A;#����o�l+��j�NcM�I�bQih�VW�k�u,�R6s	}e�f�ߋ�Il�2�Ҭ��x֓7� n@����\��[?FAkӊb���F!��9�����?y���:A�W�f�U�p��)n��Wy�K_ʱ#��sJz�,�Vl�%{/��Ï����?{������FK[d3&�J����8y�\�����O��]Xex`���3�h�j~���@�']�$k�T˺�Xj4��	��jN'���\�_�����y���O�+�/,c�#e���!���������3�>��E�V�y��{y�5W�����U�A�x��j?6ɻ��DZ	�:��/Rk�x�/>wc�tA��?���ٸ6.�
|�3w\����{N>�����M��ʽ�0���,��*~��;��Ѐz��vC���Z.��Ʉ�X^�x�_|�{8��p�e5����a�d�He�̔��i�N��JQ�c:^J�WU���qlSY�u����Q������L�Y%h��"��(�����},�$k��C���O�\`��Cxk3dtU,EK�%aiRe�vm)��pr�M��(���-�K�=�?��u]%�*�L�Ӕ]!Z)��|����S�v�z`�V61�e����	�q3����3M��1S<o��<���YՒ�Uv\�d,k�7������:v�`Mf���>���Z{=;Bb�ݼ�*�l�����ɻ(�!�����0.��9��[`���	�6��݌N��	��U�a��y~�l���Q��i��S
35�>���6'��mӪ���E_#_�j�?��sM��/�H����.�{�KX��g�=Q�%t�E�Ug��$t�.�3�l�/�ϙ3��I��n��+<��1����D�t"UY��(��
��L��Mo�-��M)�1ؗ��Z*Gw�����tkm�ݪ��9æ�����(��ml�~)�/�f�m:$aOO�
9��0T�D��~[i�:dr�J�x��<�3�����~=��
a7Q]iݮ��Wi�׸�0>��ˮ��|�����u<zt�w��2��V�0}�,�y���{�x�CsA��I+�h6������[��/��u�u��.���W_�<e�˪����SLlg}m���U������ۊ�,�����B���x������H�P֢H�A�ҁW�ҭ=J.�(�@jT�~эj�v�{�t^]�xۉE_� �����c@��Ml��G�0�c��M�Mc�4��эl����X�c��#*!8��Q��oV0�����4���#:艃�Q�|��5�å��z剪x�|œ��PJTѠ��H����̡�-�ٶ�Z�LM��Jh��ۤ��$N��6��F��Ա��ϐqm�iC�.�ڷ�z+�בT����Ҟ�>�ԡ{�+Y4�+hn���+�� ¡�Hצ�x������=t�$v�����}C�E��̟��J,��'_g`x+a(�tS�EP+ D,����KT@�.a��b�����e(APO8��a�� ���"��덞}�qT#v�F��4{�����Qi|��#�*e���1=;�b}�L��0U��2���1ݬ�m۲�cǎ��}����h���~���
�}�s����k��@��6��L����k�)X �	���T8�<Ö˟�ǿ������Ј��7���S�Y�$���C��z���h1$c�Fn�*����3\�o���g���ۜ�Y±�ئ�w�}~��J8Ew%	ٯ~��� ������Ûvc�K8�"k�:�}������uAn(�X����f㲸 +�������o�|g`|3+s��e��{���+6Q_�!c��,aM�k%1�|�\y��������~pTu(iV�8�Т�%�����<�C��X>{�����Z/1)��� T$�L>~?E���Y��1����k��j�<�������-���{X_�T]6m��-�f|�6V�>Jce��P�(�����x˦�<Mc� #�,Z��R�)o~*��tKڠ�`�Ρ����ʨ�Jq?����Y��#���s�X?�}C'�mal�5�z_�ƥC!��a�o�"�c,L��h�̞z +ZR@��}�S�D}�X��<�vK���%u����H��2Ry��-�1���4#YwM�dR*U	��R�'t�6��m��x����R����=}7Ŝ�Z#�ҷ���]�e�͜
��MZ,�j-d�(��s�v���%�8���^׃���JauOH-�^m���n�G�{�a�j	�k��HI{���˞��/n�R����k$�Zmb3!�#��-/��f�<z�ŋBjkˌ��`�9=�8咈w�gٳ�zo��T�UK���*@��Y6��KWL�S��C��jY��?����NRw�J�PkE(�5At�r�����iR	!#�H��uR�!���0��u���h����o�ck�n�C.�c��$�|T���@ݠ���\z�e8��b��[�`z�W�����B^�_��O}������P6���f��i���}�������R����͟a�x�׽�y��q3�be����ʹbg2�Ki`�w��_qߏN�7��fWB�r�F����$i##L����Wcu��g�2:���lԹ�%d���ȑ�w�K���N3v�x�~$������G��L�ʶ�	�,�	�SP[��Z*���|u7[�_�̩���+�ht�~*�[�RX[�������i���廌�y6ZvDm��%�яih�34����@'R5 ���6�ՙ#t�±u���[��:�t"p��z@F9�*K�e�����*&ey��Dv���_C+t�c+S"��긥���#��^>C�B9}�9|b�~5���>o�tÐD7�4�X<y/�ք�cp�Ōl*뵈J�e���,/�6aR��7��]$I��ȁſ�	��HM�C�[��Jlۖn�5<?�;?�����.I�+������--�e�a�Nߋηx�+�0��m�TsqJs�#_,��X�:XFK#�P�j�6�Q�D���H����и�]��S���hLx���E��q���52��Χ蛄-�n�X ���=ՙ^\gl�5[�������EO%�H𠎕5U��.l�q��g��GOL�:�X:S#��Ǫu\Z���󴫷��z�O!ZL��w=:-i������M?�4��o�y���Чp�ɖD���/�֬��W��7�ܾ����1��X��f�� +𶿺������[$#Cf�3e��	F�l^��gp���R�FsMm8� �ĩin���8r�,v��V���V�e�����@6	V�0� �{�Zi�^���t����:8�2NfL����j���.�aӈ2���$�t�ء��ٲ�{tb�����~V�nk]�,��F�[��E��3}�a֖&,I�p��pq��$j����g��ڝ��}^�T%H�ff�
|.!X�{o��9z��H���l�h
:�A��c�S��b�	5�@it���q[4'�b�6IuK�o�����g��b�W.ݤ8���M�	R�(kX��m4�/�~�1)����-�b3[V5	�@�W*�K}�)~a�4��c| C����)P���a	�\�4�ILӳ�����%x��06qj��`aηk+�94��h$)�?Motw��rd�5���u]���P�j+j<'z���)��[Ϥj�e�ѻ�g��qU����4�����z�C����jU�MZ����u���V�A�X��+Ӯ��R�j������j���u��C��/�&�Fds��o�=�yf���jZZ����Q���z�T���bq�i詣��Uc{������+���Eګgx�3��)�]BΉ��P[[S
��d��\��[�u/��E����ÑpH�"�/�Z��W��3�{6��/�u� ?i6 ��uqAV�}��7n�̗��N�2J���:�s��2�N��/�ʞK�30P �w���ezv�S�XXlR��D�vݴhw[hf���<M!�+"��'�Nc���C��:�#b�0H"�X�%�ma�#;�����J��<7E}e���m�4ՉBI�5��.9�T��yr�{���2��#�FG�4:��'d�<3�E���*g�d�v����i"�B=Q��P+zA� =����ʟ�J���L��b2�i���Bn�"ƶ^C�H0��(�Z��m�a`$>K3Gh�<���(آ���.��^N����zJ��ci�A�맩؞ԁ�%�  �${D2T��Z]wU��$���Oܧ�|tAD0�2�
v��jt���m���V�.�S�M
��O���%3�׭-�u3Zo4���y;;�T3� C�Ǆ�Z�����_���W����\��?�I����������MFG�[�xvQ1;�|�v�Ne�L7�����h��W.�jt0����*��FU���d��EXy2FK��KU��l����8bl�u�^��o��6�&hwucD�����ڂ=��\�K2���F/%����$����VFR�%��R0�kܐ�켡3}��~���j;[G�*x�R(Sȗ�1����w��-߾?��	�nR.�q�95rz�+^�3���߾ 7���l��OX�@�qY\�����S>����:��~�iRɹJ��8O�q�8�xEE��YL+�eHp0����$bR�� -M1�X����&-��,�sG�u�W�e%&t>.f~���K����N}Y���"��D�w��>E�'~]�i��`t�R���h�	ӧ]?���1Ұ�k��$�u#�V�tC�le���h�2�!�{Mo��2��Ƒ��4���)@s���ؾ�z5V"��=T��t3��3�j o�%TP=�O=�'֏ӗ׈dLyd]����
�l�u���:q�Փ���(�(���EZ����G��O��%Y��V�L�|���c8zSٓ��d�8X������E�:�[��p��G�caN�*8J�}�2NA���8�ι��g���	{���`�?�*깦�{��YYY��k�V�'a�0l��"o��=�r^��Q�s?� [��(�Dg�I.�����3�~�q�yt����W�K}��n)��r_Y%����gJ
�����C* I�8)��.�H���z����i%%�Z$g��H�hzW��D�)3(%�'E�K��bk#Ѱ�*MX	C�+ ��h�u�H�t����q��6��(d-6�N(Flvn���s�]�������*��޴%ܖ�@��������=��rG�8�C�q��V���������ŭ��턪c&�B:�.�[-4���uu��'rab4C��X�)Y�rd���:�&�F�	]�0"��lƢ�Г��c�2{�����}5���6r�:18ev_vIf�F+�-e�Ď�y�����M�fU=	�^��kF�^A���zۣ���E���	�N�@�ۊk�@ӲhH��[fx�>������J��-����jC��"a�^2�ڠ��T�I̽�H�#�d�5��~�w*��z�9�rd2��c ��+[���$����'u̜A�h��G����E��Ird26�Փ̝z���������Ʒ�uUi�uZ6Xߡox#;���s��Ӝfa�lM�A�:��Q�fh�6��x�F�n7E�M[��ʛ�
a���ZD�E�]^�)��'����:7nW��^�}��:Ϫ4T������*�R��O��A>���a�֔�`ue3�Q���i��*;,,���˲��D��W��U��\��nh+��$��|�H�'
�rh��J�6^Ҡ�ː�<¤����𾿻�Gf4��\J��;+IM�Jj��Xj|�')��E}�r�R�!��(��iҮ�(8���+ ����bn��tZ���G.W����
'[@;�D������e�숰Zro������/�������?���Ɓ�ǯ�C�?��0��������������SVPK�H��]/P�0�l:�I�G��'#�(U.I�5,��8�'���N�'Z�	@#�� ��|��R�cG�Rn�Xi�:*/EF2f�3%b���Qz�a&�j2��uWN��ܗ��_|\ˠZ�S��H/;�8���"�`[	��2q������SO�M/��?F�o�F�S�-q��B�hQ���g���*$_EW�$a�� $���R���YU���4H�}�:p5�z�>[��*���3���3E��&Y�����z���,ˍE�؊Z5t�el�e���i^m|ZT��:�v�M��@�-؄a�L��*r��o'4��|���.��Y�����[Z�H$W'��̖Б��)���Q�&C4!��"h�S[�=R! l��*Ѫhcz�N=�漄Fnl
���FN������fG*�%_��uv�h}����籲~���c��[=`�˵[�dc�|�!��
0�ݼŁk�����2K+K�r-��B�@�5�@ov�V�$���Z��7t��ܹ�W�{Pr�L
�K�QSa}r}��űdH�G�\MhDG%�j[�M]O�\���*�J��1]a<��n�X��b �'Be?�sa��C�	[���_��g(u
��Jv�s=���7������0w���l��]�@�qU\�x�����/}���&N�T��D�jtkb̕�N	}%N�Ha���]@J��v4%rJ_FAf$�T����GjH+���J+ vp�i��U�A�T���|
�"~�`e\�%$@K���= "�v�\R�j&P���HC�SC�8��i蓑�%�.KɤH���d���omV�J�%5V��iI?Q�Qc'3�WO��]��G�[�[���e�
Cx^Djڸ�A{e�o�&����d;�vȨ.&q�����Z�rH��k��i����7>�r�캘z3�X��mw2<6Au����hUBI60���h�Z2ΐBI�4�\�XB�d���#�N�C�*�)!1u�Ī$R4rnA��HEg$ ֶt:Iӵi5�
y(M'K��Q_U!#J� ��}Y*{%	laЉt���_��$��U��5��]�M2Y�N�!H�\Z�M������aN���'���MO�7���.*���b�{QQT콂bA]]+���Z�ް�
XAz�ajz�%�����}����2���dr3o�����9e�qL<w?�A��D!�AO,-�G��BM}�t555�������W�#ё�PD���Hb1� ��=/�|m����Szѻ�h��)�g_�	��`�,K�f�$�E����uX,9�H�(E�,�q���+E��$��H���7��G�����w�,���m��D�L�:B*FDo��)��Yaf&��ʂ�X&�~Ԉ��6��TRY�?X�
����d��=����MOUR)�Q�bq�ܼ`sԔ�G)��3�_A.�\�7*��T&��n�ΛY��Xl0�BQ����;�ϊ�� c�˺
����|�=ï��IH�*sMx7Z`��o)C��ۏ-�u��uqJH2���.�J^S��N��%
Q�*�p!�����h.d�t
р&M�:7]�~������C���n	<Zݙ,�/�zZ���%6w�'�L��'bPa\L+)§z�0�'m�������c3��?Z�ؒ����w�o�a��c�(��6C��L�L24�7w�a⪢���`rL���IV�(I�    IDAT]T�� A����·	�|���eu���ҹ��0�Lיy*�S�.��q������ A]�l'�B�˃b����Pk����tۮ1��|Q��i��hN�*�&�tEY��#���Gn�"$�V��lѠV��M=�|>T�@*T�'�[��Ħ-�0p�x�~,[���,��:���M���2f�:b,X�w~@�z$�Ԉ�i3�h�&,'ŽNM��.�B���
��P�����n��cEq���Nn�*�/�9ڻ�����v ��J`��P˖У9|��\�}LYs�R��ȅL8�h��Ŵr��s*��rrl��2���ߟ���P�l<V&��pP��zb0�I(�;t�R��Q?�A��C(R�T&/Y2,�#}Oᯙס�dG
�֐�'��XX�\N�޸	�AK>o�;������Rl)����H�|�����(^��!�$�$�T���G�=�NQ�G2h�����6�B�H�k�/�߫�PTPT<��M��h:`�h^��t�fce	�I;dCrX
B�zV:��bk�4��P9�0��(.di������﬙"\�q>���sE����G<��/H�J��n��|�@���4^[����ɱ�Uv��S�=Խ8-2NN��� �aIP�� {�Nn�vUD���^o�4��eP����yB���ݙE�6+/@-3V�˨��ȹaRQ�:��)*<N�NvDT����<^�d�ܑ�� u#z�\;4�਱CЧ�D6��fg�`�l'��H-�n؈����F�J$���hlm@}C֮]��W�y�t{��f��ga��3�o�`�Z|4o���"M�npD�H�Ů�ONVѶ�3w��K,�<��c��;oc���a�6�[��@P_0�l"�~ȹ�,"�I�&���edat��Rm����:4���Q�L@��,Z�py\����S�>��ዷ��r��
T��9�g���[_>�ï����2�Qt�"L$c��:0t���uG47Ԋ���s/Y��~ƆM�hh��� �'�!����=x=��[U�1�K٦˻���f[~+{,Ѱ�)E-��8�O� �~�뷶��#�CVȩJ���^#�t���tG٢������r�F�d�Ra��L��Mp�� 6����Nv#iq[Q��8����q����tQ�h㘍e�t��ySi3��Äۭ�Щ�.�ԃu>
���(���>i��9
��&�5S�<.(&l
<�,�ݡDM����J������	v,�*���%�/�h��L@C��ؗ�R�8���*��p��8��F��������핼"n�}G
����h�Ex}>XVEӐ�Z�	ǒ���v�:��\>'���	H�7݀�vh¨���q�:Bu/&�a?�=)q�9�.��IDU�yi�]��>�H�ulذ	��8R)���׵�W݄ekrx����aiUMC��������"��K2!��U����	�b�^`R��s�8����g�b���ذ�+V���I�w24�J)�.�,�Ux
y$:;�g����-���L��(���$S|Ț&\�@i�TVJ��q�iGTFN��r\Y�
CS9��
\q���?����N��l!��-���#q�1���7|�H �l\�]Ez�|��b#�Qp��iz$9�ڐd2	M�ɨ�̸�Ѝ�1��LG��4�Q�~e!Y%d

�ޥ��m�eE�]�2
�#��H�uig��p�S���A�iH�i�u㒌g
�	�2v��Hn)�/@�y������:4�_4/�L'�^/2�ǋl>&9$(�w�N�!BxQ���{,oZ����Nk��(He3��YC�?"E��" �|RZ��$�U�A@�Y�/E���a@s��0�Y��q�t�Q����T݂RPD�u4,]t-.�G���'��u�ў�k����/7�L:-L���n����މ��Zhް��Hy\t1Yr�d*�7b�Ŭ�b�S��)X(�E\+���89�(XA��m�=�=(&{�L7�և����l�J�!�Ia�ʟ�'�p{5"��BMd]B	������k����N���9|��J@m@M� t���X(^F'�<:��E$+$�!�7k$E3����1,��t{����N���!�NpD*Y5�:B
PH�k�
�k�š�C��-D<��zU7��r/^�dƀꭁ"O ���R
��=�q�yr���&��A��� ��ɱMV઻g���?�	��t�[���1�:�d��A�]�6�E]STD�Uu�hh�Wf��g����(��g!�E.t���q�v�ib�ݼy3F��{g�'�p~��B�	(!�A��n^襭Y�)|a^��[����lQf0	;�8}�7�Il>����J���?�Q�	�F�������G!���Ͳ��s�k[�$s�Ϡ��'��4������ϰ�_���n��L3�KA R/X�L�d9��?(4֜:��\� \n/ܞ Ri�o���ZE����=�*��U�y"%����J#/��pub�x܊�m`*����,8�p�zC�e	��f*2��93_�N(]���E,�*�n,�4�����~i��8K ��d�:��:����M�	�Y�H2���d�}Y�g�;���/"`�ɱ���W嘋����U#�Y �G2�E�r�$2��Ǐ]F4`�}�زN�SL�y]��n�z��-�nF*MW��U|��/�uU
Y����D"�@�	xd�&�[��%�%"�R�"��hdM�,|�!��,���b��'EE.o3��Cכ������1�l�=kp�1�pĸ�������P�P�@0���4�l�jL��A����UG�����A���I����X9m��i� �@S93��
\u�k����wop���%ۍ�~5	3�����u�~�:����h�ނ���#�+��Y��o���� kХ�AQ��w���Z�ƍ��n�)r����_$�b`n������ff+��[�nY���셲�_�"RUb�nD�.���"�7�M�d�����-�e�:	���"�!��c���4�7�nl�7�V��(���HU�v;4�U�c�J6Z&v�#�[
"?��g���c�q}p��&a*��ڐ���lm6�!����w.:�`GW`~_Q�# '3�8l2.TW�0	F #����BH�EEl�|^v1љ����(^X�@0(��%�26A�D,�@��B���~�H]PYڻ�b�{�������[����0t���b"o�D�[nI��f:�v�Q�a����ۇ�ɱ���,]z�4��Z>oIEC��DZl���E3�x�zx&����T��oX��낕�`䈡شy�bil�0Г�����U��6\h�5�B�ҝY�y����R	�P-�tN\�(���<'X� ���eV 0�v�h0$��*��N[�N��� �\�siDC>Xz]]�q��gb��Ñ�w�:B��#�M
Cӻ���*
�Ã���Ū��@���/#H�?�x<�sO:f�C��M.(��TV�V�h*��6Y�k�s���͝���z��8��c0錣��6!��+�����ie�M��_���O��>nT��I��4��y��FM!����E���E�dd(Ru��TqW��p!�ܔ��%�4j*��h�.�ӊ&�ϫѓX��]��nE6,Y�A,i,�/��p��y��ƛ����O>q3B>`�ǝr!�k�9��Y�uCXɚ�:�л.*kӝ��Ӱ�u����|��� �*�,��D��ۯ��5��Kr�⚛P(�)F�g 9
�y�^С��(�N,6�q)�ln�Gk��X��rtu&�S��J��±�D/�K�$`�����q���8
c=#A��t�(pm�BN�6}^��z�|;0�9/�t�"�ZD�B�<�T̞�"�;�x�u�Ltv���^WՌΎ6h>�}����#����X7��W_~!�����.^��6��� �ѥ���4�����`��'�����"�^�B;%�:��ɘ���t^W�T'<n�ׂU���t!�MK�j \�d����@��Xp�1�蓯��_
�f��@ڬ-j>wڴW�	�6�hk_tG�O����T6����N��B��fYh��#�95�|,]2�=W]vV�����B.���o������ޭ����K�M�f���L��j��oHR���H$q�G�4n��mrA���@S9�����{��yo�Q��=�~�l?�V�[4"���3y�Y��/�н���њ(��͝q� ��y&>�d![�#�+H�*�=�أ�Rw�����Ի"���ۮ�)��З�^fb��l;*�-��.;�ʏ��KU|i<��4D��Y��+����D�2�{`�0�xN�t֯߀��8C��?�7?����dg'��-�4��B"��B�qA�Z{<��w�G����<��Ǹ��+�Ӽϱ����'�E{W�lG�W\1�hR}�7�2M�Qd\PT���!�FW�fd��ѷ� �j�o�lY�뮻{�5���N��D�����(��,�T�a
���Q�p���)���ȟy���vjxB��ĺ�ϧ�&9�\S�QW��׃������A4T/mһ�:˖��}����nJ�Q��מ��3�F�.�K��	��	��Ew��=z{\0�n�sߓ���wF���I� +���ȱ�i!���%������Dg2~�D�4L�uR��d�q���i��:SQq�bm�l�4�"�оe#����3���۟,�M���D A>�C&��b��Q	��/2w��a�S ���d���d����;�L:��I��׊y|*�;���8�1�a�b�ѰԐ,[�Rr�ڶt��:���c��!p�>�|n��Q���g�m�E��)
�a��WD���r\�9��Ce��
\{�����ټ7u+������Ы>��C$���5k���O�Q0
4pV�X���F< �|^�o��f�5�-#�3]b�&��}�x�$c��hش,��&���H���FN%v��f^�����S��S&� ���t_s��y8�m�ƃӯ�ϫaC{
'�q.F��t ֮\�'��'t1p�Pq�!���E����O?|���F]0�W^~;���S�ë��+s���v�cot�^���&|�+7#��&\=e"�<0��9�k�L\x���u�^x�ݏ���>�+�H��_|�/�Z�p�
�5�< 9�I�X��55�xt�,|;o>�����h:\�Fm�6	��Սw�yO��P4����%Ar���aذ��F"������8�c��c|�N8�D��݈�7H���o~
 -�Ą	砵W_|���X��g�cX�v%w^��3&��co\}�Y��1��o�"����Ͽ�/?,>���(���b,X�����ك��?Vl�׏u��$$q��UX�n4������w�][22����rʍ��՝���8��E����Q�҄x2�ؖn�Y�J�At�e��J�Y�����:b^y�������:�]Ix\�6�p�ֹ�!��R��1���Ν)W;��� ^�z욃2 ���!�H7VVx���؄=w��/=	�\;Z{a˖�"X�o�%uo��6�v��X��2.o ������
�_����sN9j����mq=����@S9/��
�x�+�����7ӹ�^f=p�x��8�4�a����L���h��d<����i{tvlA�r��W����pox�ER�6օ#��E�l.�Uo���f��[�h$,�we�����љ��xE�l�՗���R���;�@���7�ƹ����?D"�?��{\�t<��hmѐL��v�U�s��o��,^���4c���_k5�N�nEC�Fٸ�S<��g�������b*�KA^��+�э��w+�4FE�2��+�=���@���2x�gз_v�q$�������t�l���x�;1l`=��X��b�����;�yG Ō�n���^|��2����0�u�1�+W&p�q'�+.���탍����R��x�1�~�ԁ<�BZv�a��:�6�g<��#h�U�S�8YFP�[�}Z�Ϙ]ѯ_��[���_��o����B[w�S��_.��;��~+�������5���g�y.j<��?7n���6Dkj1rh�)����Y�<���{�hB���e�hm�u�x���1gο1f�0a��H�R�{.o �Ia�tvq�}O���_�{��;�����ށ��ۀhm_�Ae�9D�QXV20���lIs��$"QR��%��
#�C�[9��,\�s��gbm�ӄG)�=��q���#�'6!��+��� � ~Y��*�M��n�vP&T�nK����@*�FUC\>����>�/8�R}�M.�����
T M���&+p���������&r�����(f��S��ݫ�֭�������$��:\���f�5�c�j�Z�M�b�u���܅�n������
MKy1� <�2�R,[�O���������Ŀe���W�7{�ұu�q�D�s?|��[xt�s�e��1��X��W�?�f�2��T���Y�i�R<��܃��K0��+�����o`6�K�)�b�����x����ԈXG�_~9N=�$��Ȥ�ۦ��_���>(�ҵ�Wtun��Cj0�k�u��}�}4&M��	g��\��g^����Q$c]��Λp�Ac��}���p��w����}�G�?�77�~��+��3fw7��N�8*��l��gM��e+��{���B��..�<�/�#wVW�p�r���z�y�<r�=FBؔ�;i"6������i�&KwV�F&\�T��*?v�m477#�Ս��7Æ���mٚn�v�i�����p��W��S�����Fdb�8��q���#��b�Kp�7㉧�~���&L�z��X��c��=3�@����`ƽ3�ȣ�D'���2�J�[�3N=�H\y�Y�����/�
gZ�AU��2�Z��W�{��w�^Gx�����;��w��%�e��0���ѝ@��x�l`��1^�N�6.CĿ���*�E;j���T?(N� ���N.�]��5c[��{�,�P�E,��'�|�_q�����EO�v�:�B�Z�7�x��>��g4�*�8����-I�u�Ћ!i�v�h�:��]/<|�w��R9He�`*��rZl�����{y���k�h[�7\>��|?�S��Ԣ'у��~���:�{bRP�Ie��;���	9�B���;u�:�!��lr.��#!e���L���Y���G(�ʔ�hD��?M�����X�YD"֎}�0��"��?� �{����x��OD��нwBѓ�F�8�ĉ�� ��r�0��|+W�Í7]�̛�W^y��}z�6�;�AM���1���x��i��#��p�E�a�&ѪSh�J8���U���Cp�C��O>ä˦��xcGm�S�E�>��\
���n��2�}�I���۱j�j̺�NԄ���s�U��3G�G�G��ݷ��x�ŗ^�C�by�0�oG9��r��.<��CP\*��n�I�MD(\�����Q#1���0���Տ���G�v�����c�'����w����L��;������Ŕ[ے�
c��a�=3�д�Ϟ�(��Wݎ�oDU]�6��i'��9BZW]s�4�_s��Hf��3<�0�\�y ���a*��/�\��_w!r&��1�����.�x�=z�8՟}�C̸{&n�v�ta55�K֍�
fV\H�θ�E,��{<5k��x������	�JI��OIQAw���%%;�Kjp�OFg�5v� 9�iߦ�[��l@.��)0;Hѥp\E7�/�վ{��7_v<����h߄�6�𣪶	_�[�t&�Pȍ!�`�w,�"*�槕�t�P��j��;O�S� �mr5���Z�
����dn|�߇�<�7��nݯѻ�{�l�Ǿ    IDAT�BW�z	p[��.�DB0��?	��hh��^���k���;D��,���3R���{����"���%���h��s�_
$�þ�k�,]T�ˁT�c���]y:�.��<����H�|��"��3.�rCp��у�O;7�x=;`'��&&]|v�u7�s�1R�9����cOëh3z7\u��0��Sob��O1��;�����qٵw�i���be57,�w]7���C�*���w�������O�WTCۖ�\�(�._�>�̼�&�Wy��݅�Ͼ@r{^|t&n���;\y��6� ����q,�>}��t`KW'V��FK�aX�|���>7�q��Νp<>'�~�c�|���3k�/��)��ģG��>�������`��{���}���<L��Q��^w�����?�9s� t�sNǡ�Ɖn����}�����CZ�֝��SoDWNC"�����O>���*�A�ǟ��Əǉ'�C� ����}�ST�|8���#�����܎�������.��a��|>�����+/��a�(��8��K0|�p\s���f���~󿚏ƪΟx�k���r��+��λ���G#�)��g�¬��Du� $Һ�cZ.��!�bIB!d�4쎰S� ��m�y]��I[;�L%
�E�.�v؞��L�v�Ȧe��K%�9�xx�dx�1�v��uk\�w%@׭۶m�f��ضm��vlg';�m'۹�����8����ZUs>k�Q�S!�O�'Y��/�8vE�w�k/ż�b�t��6JWU᷁e�+	�d�&t��)�AWV��U�.����%��|�YBW��D�-�P�y_��~6!XF�&���X4?TIW7�<r2����ۙs�v�S�GD��K����
���FѸ�3Z��^�J�e.�r�Hha�qD+S(n���Y�I�'��xY�)�M��'W�������wn���7�M���Z�j$���8Ӧ������4=3@�"��Pn���E�n��^Z`�NU����T� �$�ڔ������˽7^i	(����y���s��%���a���ͭ(������C��~>oG��Ĥ�8�������K��!
�_�_x��d	��)���a�wB( ��������r���U�p�\rz}�?Z�ܴ�I3C]ԃ��n'(y&7k��L��] �w���;��d�ɭVۃ|���ۓs��7^����'�I�}�+5Q,�>�R�^Ht�~�����=*�u8���v�Z�8W*�/��s�����n0���߹6� ߫v8��hEە��?�@D�0Pq��e�,�9�,�o�E)����j�!gg���_�!N-�>��M���s9SyL��=�E��1{wK3H�eX���+a��XY�q�rJ���$tƳ��
��G�W�D^7�~_�̳ň2��j{�Ͽ��F~T2�m.�Dv�]�y*�z8AP^>u�'�h��s��6��d&��Xg'О)��WU�;��y����x���=�(��|Y��*ꭅdt�D�o|�F�J��}�`����1~J�����E[�-xC#�=X�ҍ���m��L]�KB/��zB�w�&HU��W�p�D��`����aQŠ>0����b_�3vװ�%-�`�ĥ�%C&��m�R-%iu��)�ɧQ�U!T�8<PK_um�����4O%����[`��h�eW!�6��:	3�ܐx�X��!������5�/� � ��i?�����rð
(�FP�|Oħ�o�M�K��s�+s_�>��d��ܼvh�[T�h�׸�B�Q[���������"#�t/|�J��84�Ar���\��	�I��I�����e^`�5�w^RA�@9������:�. �֡����y�KCb�/�o��~�f� 8��j�� �;y:x�~3��i�z����]���ӓ��o"�}/>��HI=	:s;*�A� t�RE8I��t�}��2�x�%��ob��\*�G�ʖ���l�6����#��a%PÄ��?mĵ�py�6�Q��n�LnO�^���;E��&#��N���'B/��z�@��Ϣ��O$E�D�ۋ�ky_dN�ݰ�gIq������[��Ma��n�#�^;(UZt���x������^?�2βg�1%O��)؜��9e������=r���	�JK 9�p̺�z9�Z�v�'� Ե�e������_ �Z� ���Ͳ���#��=q���CƦ�j���r`������FӶ�D!�L����;K���+)�>l�b�QK)�<F�C��jl��(��É���1eI|9�V0a�� �О~��H��{�RV�� �pF�k��i�A��Is7��@�d���SL4�j��-���,g��T�:H����$���l��q�d�݃�{��6p~� "(_���pv�,�EǸ����8i����[�l����%*�#�O��u�8��1��?���P%@4H2�F*������%����2��&���z_.�'����B���=�`��\�^��d��v���܋�� ���N��Ҧ+yit��9�N�NL��.{F��{N�J}a��ݽI�ee�V�"�Q�߭���<��B�+}�;�a�h=�-&�j3�sJ������J��(	$�'���?��Cz����=�E8���h���q>>+7T���+/�&�x=��$�=�+�B��/�f�^���O�Qs4<� ��3Q�����%�Ydp�0a������_���	��(q��ȱ-����r�*J�T��\������lI���#��ރ��A���� X���:�n~�$����`|��7&�T��<?DF��s ;mׂAw=����䌽Pء���q��[�E"}]{v�_'����u;jW��$0���U���gDXhb�������& �����ـ+���ex��T_i5��Īl��4�}�M�4&�X���U���x*8:d%�B�&Ѣ��<ڝW��Jo��勤5s�SϴHl�2Pc�r2ܽ�듖�|�����~p�%;�kSbW��(�Җ�C"�r�=�z�ܛp��76c��C�&��i�PBH��5^�=x|�5�6����[(�=/&jt^�!��jA��}���]���O�{�a�zlSlY�[vܞ	�i���X��d$X��p�r�"�Vle=x�/����Z�҇X`jۊ %�F�r"�ק���:2�x��M�uk�Z8�Y�~;`�>i�݃�V���g��0����"�I_���j�y|E�	RP0g�v��g�ל��ӏ���K`�+�2�3�	q�R�l>�<ԽC�a���E�,�\N��Vo��Xh:��		�	�'
Fd������!��Kh;ff��	�il�<��ia Zg|9����#�M�;����i��H�+�����$�25}�z\�L5Q�j��Bi9|�^<�*hDwN63��/X�s���7���N7B�I���L�����X,Y��"�� 
.�M��Pd!����/db!U�m�O���F^�;7��߫��_�Ȋ����֩V�̆��k��+���������������㒖�����q<����v�&�k��P*����͔M����#"N�_~����FP�6\�9:�X^�o����ME�/�|)��U�� Čyv㡚��\
�P���'O����4j:��˽�<_�v&5�^l�`$h�E
�zhzQ�ԟ!�\���W��MB$��.�
2Yf��ul�8�Z�!~Z�y�	��Й�>������'��������lZr�0냵ʺ�b}�5��CG�������/��+��3�Y��O����~����0V�8$T�-<N�k��ސ>vt/֜F,�2x�"�� �Ưs'���r��sH�#�k5:tدo�j�Vt��]���b0h��E�Y#K�Z�Z�H���	(qރ�a����n4�����4ʾ8)`�G]B�!�Ғg(�?�Q�(�|SY�bZ�a�y�����T�2UT�4���Z�i��\U�	�R�tO�g��;9�4�����(Sd_���`����|�g�ڿγ}^���!�$��h�Pi`�!��w�C�u�K�Uw��^\�>Yl��o��8M+V��%U	�%��	��V��g?��u�~<���<4��2����y�����5�5�=��'����i��/��$��0�����\����x�@	�hח�x �����u｠�iO���t��;��f�@��\�.��Oyؗ`��>�Ż���"C@��Ŏ��0����:i���ڜ�W6��"~�(����J{[6#��4-تNO�-Cv`���4Z�[���v��� �2g��\���"8�򏂨�1���:uc4Q�L$��mU�]���q)[�0,6h�y�C�{��M�G�Z*�����84�&vڸ(�4�2(G��IN5@�݀�x*�g���� �
�'o$�g���d�V�'�$M�y�Bc�G�=�|�7O�v����\��׋�l�Wx�4W�|����E�]f��N�6�����e5���"���E`l|Ճ1��=�0Ax�]��v�d+�ƾ�Y�����>a������1	�����J�����B%�:_�D����ǂG+Y���C祉�CE�=I�s2w���4W`��&Q&rL�Y��.�!��8���l�5�p<~���Д���&--�OXj�����xf�䨱2^�I�E�%X|T$-�\^0���8��f��5|�nҺ�t��v��z�/#x,�F�Ls��2��9���0�k�s۔9�3�����"X�"d�rhL;���~���z �~�_�!����p��v,���A�.�n�!�>|(T)m5�B�]?~��d��I��5h
��y�գ�4��N������A(�t7��C�����a�,R(@!7�w-�0���d��QMK;A�M��,�Ɍ�P�H����Ɗ��h�7�#�C���k��l���: \��%^�eM�wPi)[9'�*N"�֣�M`��#D��Lݠu ��ѱ3�}��o������O��P�������-��܈�@戱K)�E��}�y���6��d�*8/���Z��0�e��2}g�퍙]�z���1<�����N�-��1������^3���՘���kjk�5��A�Yݔ��M|�y��ʸ�'ļ�M_��۫��q�U���/�h|v����������,��:�Z�-/Tܹ�Ę��?���Oa�	x^�%ڟ�lf�@W����&Q�3��57܈��ؘWݮz����7D[s�����?R�7�$�xz� u�׬N���Ӎ� �u���I�j��8�8�pt���7�C�z;_\�4>?�'��B���t�@d�� Pp��W��j���>>��*CȽԕfRR����h�!(F���Wp�wՈ���H���*a=z�_~BX>)��N�0�Lh�N����66�����u�=.:�%�m+�%|	�0��e�;��(�\AAaG���7W.$�	�@i�36s�H�@�">w:�=����/st\U�/J���RvY\�� ��%r��h�8^4�QY|���i� Q���c�Aڰ����JY���-�s˃�lڡ�cMCd��5��-<𵩖5�@S�p`V}:ؾLk��[8�;�Z;�.k-�ߚ��D��@2��s�|���A_;���&<�����F�1�kw� ��~���.��,�>�|J_N������z�,|q�� �<��=i�60?��WǞ��#���Q����1WGlM]�،�k��3;4����Sݱ��,���LD;����]��
I�Eq�N�2���̆�[/)�M�_+�~�:�v������+S�aE�͐���Z���>����)3�B�ނ��_�Wv?�g2�?.�f���ф�Z���}��6����qץG�,)�_�mm�9������oY��Ւ���n��-σ��mp�!L-���d��Q=܁�00ќ1k�2�5����FE��Ӣ�b+���*:�X�����1*�J,(����I#U(^� � ����S�jXJe��6d�L�`�NM��{���nI�H�"�w-l��D�9v�D�w=$ NdVf���T|ɍ��'V��i�áx�	+�ӟ`%R�!�;%�uB�v���dŲ˓ؑBo���`sw16s:j�!ܙ����1�E�YX�\P�(9�է<Fk ب9�����v��;��c�9m�/\����:(���ϟ���=�us����l��7�w���iL�7Q[b�X�/�dͅ���W�d�2pk��-�+a��Kw_�'6f��X����˞g���^פ�;,C�O���L*d�4�?��7�~�M�q)3�er.j����*hk��$��،v!����M��Bɧ�a�LAC�^F�2D�(�0�s�s-��>v&���X)�OE	�&h�Ƅ���ڕ1�PF��p�׆܋b�E�@��9����P6�Ae����J��:C�0 ���MK�N#'�h���2y�m�3�õo�i#Q�g�!��ϟ�����x{��U���0 �6$F�g��gq���"40�{�w�9��/j�u%o�HУ�pԢbc7�.T���x�L�\1���="N��̏**�Ml�Υ�L�I�>5y����4�j�oq� 0��B#)S��%��ܕW�tU��\��=u6���æ8`P͍P����OX����/؆y��V����:�Úܡ��C�A��%��KF���gQ�2$����>���If�4�:�h��L%P+)��lR�(���!����/2Z'��"�\.^U�CĬ�O�PVxؤ�~��5N�6���$�Fi����v�'XG��]H%:,uf�58���=x��:��c+�V�3@�;��\�ds-��J��Vؾr�m-K2VF0�.�#9=/��4�U<a+��/7Ax9��G��Q��f�vs�=]ɗ(2���
HH�����͚�j�#GA%Fj����5ⰰɥ{T�D�������Q!>y�����i�CRf�n�>h5�V���):��,ʳ'��"�8N�iM#��M�4���g$Vs�`��0����>���9u���N|��Q�nm6"6EpN�����S�aTE"�Gu�Ȱ�Q��0�����������?Ը����1�~�T`��a8����e)�Q�A�$�\%V;g(&����,�����u�3��ŏ�\�t?�~�w��-�\��Uƨ!GA")��!Ϝ}(h&UC����	�Јݿ�.:''���(��0�o�xs�|l��ú�F}���˯���C���}�J6e�D�^��8t���nO���@�ת,�$J@�!Wd��� fl6/���g��u:������&�x���W�ׂMv��M�gV�|S�ϑ�e�kZ�f����!�&(��ww�:Y+�x�J������D��aȿ���VrV�G�?��޼������Ǌ+�j��'?]m�C2c��!t�����`����T�Mr���Ny
�|a@R´i��-�j�������_R_��� 
���)�<SG�,�kv'ُ݂�%px[��	��ư�ړ��iT�T�^���T�%ؘ��#�v�(A�� 5̈́e��6��
D5�&��I:+��8�*��M1��y�{�!�U'�G ��h�)Tc�_����d-���=��ج�m d����/�@B����)�j��Z����0�-�-vߒQM4�E����l@�r�XB�|
*��X�%4�L���0ʡ-z)@�~����
e����\���(8�Jcx�7'-�X/0��$�uC�%�6��n�(Q�1�3B��)�Б���~�{wn��u������أn�/��
R�z�@2ICk��D��c��ƍ��
"�/���.�N�b��χ&R���w�Z� D�\ޑl�Y��';��,8�Y?W�G�*kl����ˋ�8T^T�<��wxgoe�ＡԵ$!��W�!w�%QA�bsG��%Fl\D8�F$A��?�ܮ^�f�f?�7X�_�d�Oσ��U��f�$c�q x��	�ިʆ1��Y ��Up��/_�uz�������.6�7G+����g2G����,�!L�����߲:L/���7��ק���؉�R��z�ճ����"��|�}����T�T� �ՐM^WW6�w�&Qc���ߤ#�<�-�?��k��}�6=�����"��9)����P�7* �@4~DI����x�Rb8�x�m�7�����	7�4*(�k�/A�O��(��1���#6ݵ������`�"�7�V."�51���6Wf����ot�4�e8X5R����^����FC$��T�Pz����q-[2�ht�ɛD�
>���P���Aƈ���'w�}�wh9[6j�Ld���@W���r���L�J�+�_k���/�F�ϐ�_�]Ǿ�^y�&�+��]:?)Vo_?��1@������;w�UIQUC#*������V*����6	Y� -��g	q�� %p��_5/'��Vm`z�^�d0�%L��/�{e�K�:E�T�s��F�B}�����z���u]�����!Ae.H:�""��#�D�PU�,����F��{�#����5�ֹl�щߪVgK���"\y��߱uR�7Đ��2�0L��b��������%�op��Ѯ���S�4"��XK�I�~B����X����eڅWX6ٹc7�[�mi���+�'d���X��q�8��Jܧ8*�~8�(f<�U2 6�̑ۙl�?s�J�c��f�<�--ƻA��*_���7-�K\d�r@��3	�g,	2�t�$�$�,<g�t��F��A(^���y�Z6SU����@���s�fp5��2��'��OW�#�~��ŽR̍E�,�j�o�z��ěq|>q����j�u=o{����	9���ǂ�_V��m�*���Hm;�Z�΍��?^�n?e}�>m���[ZS(���Bԛ5����4��>Ğ��~|��3�R~��9p5����<��ڡH'�0Ef�I�YoP��M�D��Q���ȃ�
�%�M����������?�f�"k�Pt���8�a��r8��p���[z����P�쑪�#��Y_ײp.��l��+[�Q�t�iۄ=����x��D�Y����Ei3p'J���B�`�V�.s�x�!���*�eu�'��C�yh%o�w/T�u ��ߢ���4:#�&��J�����J�`ӥ��1B^�NLF�E��G���Ĉ�2��8`0�l?c��¤�Qz�a
��MĞ>]\�
��"ʖ���Z��ӭ����z��l�6���U;Ƌ�x�)��x^�5#�K7lT�
���%��[�/��N��R^�����/T:���\���0D<�$8��SGMM*ɴX��Y�\A���q�z`�8,��M�_�ܾ������A�3���1㭏r歑��9S�gN�$zT}��NM���M�A���O�6�+X�~�n��.�kN�%���>��*Ɖd���w�t��/�i�z�����i�<F"��h�E��P����{>�<y�Q�����b�>�|�cL_-S� �ډ��O�W�[��@����O��a&t��B���p�S>��VaZ�����w@����ˋ�i�|���3F����v�|��-3��<(}+��&�������	ƉH�ӣ����}?#��T�l�
���}���?&��&���nIS?U�u�MKmdև���j��"��z���|[��ȉ�Uѷj��*�/�
��(K��]�� ����j_TF�uNH����3���q�
#S��˿К�c�$S����K+2ݯobu�
���߸��u�S���J��&�qDĂ��M�-�J�*F�c��
����� ɻ�*�V������4���GTܟq��SN&ǜWYc)�l;4��2�4<wو�@��L��2h�"�b�	�8�%�vg9?��`Xg9�%5�D9+?�"�Vv*ڮN�]eƬ+��/5כ �qU�����%fK���o���qu2�9;'��(�E�1	Ѫ��C@HZ�B�A��.�XǳlW��跤�����T���r`bq ◙�6��<�#��2gvQ=<?�Ǧ˂��i���M�I�H��_��>�R���Li��M�oN�wF���� b��t@�i���!���gn����Z�]�Q"#+�)�T|�'�:�DITL	�o,�0g���#:�&�d�[�e��D��ֳ ;�s�����AΧ%d&�e���G�}�Re�L���&�U����P�5b�Ci	�^?^!�/JUY4��~�U$���ښ?7��FV�Q����DX	u�=p��Y+(��>�qۦl%D:jC����%¡����QF<��
��;��]G?�G=�Dgk��V�}�^{�׈�\m*ڽ��o�p�] ��<ܟK*d���J�!}�#�QɃ�2��EP��뺷���?�@~���}(���h��^«������
�����1���a4�8��g��C8pi���s�%����y*m���ZЌ�HеBX����b��o����m6��?*V3%��V�ՓSb�U�����Z�D��7�?�;/~e�K�o(�k��ݽ�?P����ҨЕ��[�6Z=HЖ�>ݛX�Ag����ة�!�����u�I�"A��ɚ	��,�ppU]cج#��wIZ�@���eM�+��m#aXx��j�v�(�l��Y�`�L��P�Y�P���x�3f�2�����'Z �3^/�@�f�~�������j�p�C[��#5	��v٥&���T�&c&�o�"�����1�mm
)��(�8�=��b�G�t8 �;�Rޣ� ��mL�=���u��f=�߽�x�/~&��K�8zBc����;g����)�oQAb3���?�4$��a�*���� }n�h�V�[����K~���F�ђ�W��m�kd���"s�q�g�7��2�	!h�",�"���M��3�#�U-���6�$;-`�"j]Lp�:��;~�Mԣ=s���թF��
������{��a��K�&\����P�Q	��1��[K���5�Ė�7�8�.�N��Q�Ó���&)n���)�Q9��|�2����4$z���A�6=���P$��:����YyE�a����RH�
��0(�Ƕ�έH�� oPM��:}}o_OIPHX�y��Gah�-c��ƚHx �R»�v�T�ϋ��-� ��,�;�Bh�:��^\_V�2I1�А��� ����vU0ybP���V�@�[��"#�u�譪��Р�p���"�Z�_D�ǽ��0a�^�H��c�����1��]�rd0�#vb���y��
�_@x��aP$���]c*"�3�RA�7�k���R�ReJ�F�*�y�m8�SA�ߐ#B�I���8���>��%!�*�L�~yy8;�>X�$�2X@�a��w�V�� �����,�d��M�ʼ�����������@�Z3ެbG�-S��<\Y�c-m:���b�z�oC��J*�/���8WvoȟK�p��pX�x4���g�(��=A[�C#24G�Þ����(�6]�z_}0�rB��Q�,���U���ߋ�/�{�cT�@Y9�"�Q��s����?U�ۆ�~�"_��8m�W�H��^�r,o�������Lh�ӊi�U[���6O�f���U'[�k��~����Ǐ{�ݤ`lL1�����I�����'}SBL�g��1l ��>c��1~{qնn�kw;Wd42<%��iؓb�j�~{�URi�!M1DS%�g��9k'���4��y�4�(��������54�|�Z8�NS��[>�����~`^iȚ� �1����"�FG��1��]Xxxa���;�l�bY���c�R�0f��	t� A#�>��"�[��}p�4)pc��D����L��$��~I�<]�\�+�$P4�2��@�g�y����h��`��4���'\�#Z�68q���e��]��	�{�Tü�`v��j���ۛ��:�t�W�ꓠ��O�+?S���/Y��u�1
"V�fF�AS����Cʈ���!��D�N(��Aʴf����Q�k�.ɂPd�5��"��}�bB���+7!T����`��t
�Ys����眰��оoL"�SV�xO��ɉ���/���g����Ƚ�X�hu���^�<

�\�51$J�P��Z&/QƧW���c�\�4�u++��1a˃y���0�2ECau���m���wd�����v�/�/��ȉ� 9�z9���	I:�/X�0�!�6Z1��|�L+�~iぁ�_{���
�FE��:�b���;���Qj��~r�t�ӘU�;�M:�2��;����=�ڿ5_�݈���D�&�D�$�Q-3 h$P��L8��ڏ��+�:�D	����0p��oe���$� �(`u�s�*	��f)�|��y���{WY~0� �E�OG�GC��+M����Lz���L%"PM�����
;�l��=G���p3aTb�9�2.�I.w|�����Ru�R6������� v��g�A�t�$���!��XL�^k��>{LF�L�j�H��]k�[�j$��Ix�ޡ޸U���x��}=Ս�n��/!~0Q�5h�/�R��۝�o>�)tV�P�ـ��]_
���PD"s��%[�!.?&�tLv�e�d��DJ���i���ԯ�,R:�]T}I-���H�H<��A� �52��9T�ˣ��<�v����~!f�/��=�8}I���2s���މ�L�}X��?�9�:ϼ]D>��^�5���"�(c�/"eՆ*����+k��z%�ҥm?����⧀���X�N��,��G��fk��q�w���&*������� U~){�^[H��2���v��?�y�˔ؿ̠�Y�ܦ�W;��\ v[ݨ4kVYKp@��[�AR�ױ�MD��Wɣ���P���
q����-�7ju��Z�(_�ޥ��)Pz�8V���\(�IW;!�Oa���d9
�r:L���Q�7)���T�G�j��8)S�cVMu��噽	"ݘ��^T��ԡ�)����Q$9O^q�UDv��J_�e~p�ЊŃZ&HV���	�^�]�����[��X��Q�6�cs���T$qV��P��QW��*-H|MZ�l��N�b�a3��r2�L�����=�]Ee����=癯���D<�^�z/mC��m�i˹9���`H��'��ND��!�":l��?B0�8�	V��{-L���aCw�JK\��ŮȾ!��91:ڇ�qg���BT4$���э��L�w� ���[H�Bљ)���e=zl�A���c<�e�x~89>��/�h���+Af��2���&� ��Sw�U�)vkۡ�����_5���������e����=�Z�b��af>���vR��\�\<n(�=Ycΐ�Ǳ�O��G��{"�l@L���k�f��8�k`$�Qj��}�B|Y|�{Y$�mX���ؙ�?��w���Em�o��9Z&Lڪ���������*���Y��npDV�-�eӝ�������&|��=?A5z%�b{����؄+0�XH�}VV�^��(Py���q&^�%�Il���;U9��kO�nؒNQj�$�]��y����0n""��$� :��z�v�~���a~'u/���C2/��x��vӱ�[�%ִy���"5�e�()��cV���Q���[��2�"�G+���|!(���y�x_�I=�MN�mK��J��4��hL���:+���K�-E>ӢC������Ƿ��P�֯�R<��B9���:�5,�8�u�~��1�B}��Q6vԘ�G�%>8ہ!hn&��]>�h��Zm��и*�����5�ǃ�r /��/����
�J��s���ƈ�Q�(���܅�Oz��F&�7?h�w4�â��D�ä�@{��&�T����n�g"%�!�>]� �ARB���e�,AH`c&~��GDA_��J��{1'�'Du���د�|i�/5��=�ߜh�[z­ҫV�AP��l{b�+�d>�Ŗ"|}^鮚^85�4�?l�(��ӂh-�ޯ�{]��8±bD���T܏��m�:r����j���[��|<MRN���o�P��fu�(빿Z;M�b����@V��Al��¨�/���{�	z�o)��#IS]�b؄�ֿDox&���,MU�����٠V�ù�����*B�c�*0,��[,wД�o2KE"�k��	���	�⽥��b*4�a���%�6�ò����eO�PX��g8G3n��ʚ��ﻲ(�C�x��P^)U9��G���H�e F���$�Ö郵3�F�fďD
���
�ǟ���D��˭��R�(ʸĽ태(�� ��#}��q^Q^�`B~� �s.�1�op�?.�,a*0~�ȱm2�<�IF�o�V�r6D��ye��j�NO���+꒤-e��&(P~����b��?���q
R�3�V ����J8��р�>�Sub��,�,ƈWf�D"��^A0C����/���	j�sM��8wr<�9[���)(R��s_h��iJ��g\^��UK������[�-���x���a@u�i��Z�+\w���ԯ�~E�d���N?�	/�6/&�^�����Aǂ4���(h�9�L�t�\Wz�#s{P0���LEo�b`6$@k�(3W��m��f��6eS+��sX����bb��c���)3&��o>�n�(yfHО8������`��ȴ��%��?���ab�p#�\jQ��H��D:������`e7f=��J*h�R�Tt���B����-!�ȊnJ�������"��2�=��f�l@�3���Y�I��'� ���� �� h�I���V3��� ��I'U�d�D�d�8�ߛ'~b㽔H��f�O�6��Y���t�:
��������)�e�(��x��ϲ9z�R҆p��Å�y�[����),`sr	���`@}i����m�eL=7�78O��HC��4�2��F腢z1�|[2�<urR+�#��4��MI��ֿI��t��CĈ��&�e��`��rr���y��|���Pg�~5i�pD�2ZbB�{���\g�Y)}��b'ʟ�E�;��UΨ�[<+!��z���1Ɨ��s�	R�~��/?��V���%��>^g+bC�e4�=+��>��8�G��~C�Ǯ�������u��y;R^0r�(���e��V��*�@��%�����徥�u_@l4�� ���/	��W-�	�����,fyq/�CE)�?��WVôMx��
&��F7��dP~�@H���a�x;���o�(�zlfӴ{ ^�cf5��:��pZ*Y�W���*�Pl���I�Ȫ�n˱��?j�]���v�AzN�02�x/�N�,���p���� ]��@g�VLsgIUV�7�@{D��Ǵ��0�[N�Ј�Ǜ�+�!abY��`�A]9����q3 l�^�W=q�D���T����,���,%���t�&���FM�3��b*���}]�z���찡Qf�P��I*M�A7�˫%1��01���n��V��+Ύ:/l��H�yT�mZ�m3�<&R��_���W��Ƙ>��*^L�Ͽ`w`%s���(K3Ehu�$�Z��x�H��?a��%.�t� �o��zT���J�\w����^�Z��o�U��!]�����7'����;�q�.�o��G�(J
%̬�@���r����%���߼�Ɗq",=K��V����R��Ҡ�����D�E����Q
�E�k-Q�ڐ��c��UyV���F�@d`8"���U��睻+"lM��=���ƞ-L�R_$j���>"V�l�������\a���5%	o�D�_�`I��q��@�g[&�4r8_�F���j��G�>�T!S(���Gd�C�X�4B�SVt����d�Ub�6��e�L]u�,&���Bڐ��k4�j-�1�=%z�}����erUi��ԙ%ݏ(���HӺ�y�98e@���W��t���cД�'Nc>��FhD�:'�����D�/1�����, /���h#t9KP�)��ɀaS�s=��f���@]l�ȵ��qm�#�;�h �k���\�㬀�~V���T�T(ܟ:~�Z'���QtA�Z��}'?��U��qz��M���0�'�ݚ�HdY�^!�((!HN2�
<CP�+��J����kW"�o_�%�ŭ=NM�;��8�<��I	����cgAFM�צ�Q�'̎z���߶�M�!Mu�y�o�Ւ8~�����ϰpu9��=mɰ<�_��ؕk����JB�Z�h�F��`���R�K���u2�>d�!Yh2Ҙ���~5�2���XС���N0I1��� �;0vI �!B~
{+(w#?J,�����ڄ_V8c�ә�3t6$��@���=$w'�/���ON_O�p/^��
*��Й;�Mj�8�_K��
>�`@5JR�����刺`��n��

+Y#�H��ň��������T�]\`HS����|=�E(,�3�V�J �LÆ�`u4�:�D{B�f$�ߊ'Uj2%⚼ԑ8�����w��?jY9���3��?v/���[p�9�"�`���pY��T�@�N�V\���/ ��I/Z��K_h��R�ghM��$C��]�:�&�3T�����Cߍ�3���lo�}X
�=�@��-�W�H��z�h��:�����-���"4E�Y�vC+��C L�fd
uq%i0�N@(�A�P�A�)�($������}�k���������L7��v��?�*/z��F�\.w9��)�����	�t#�i��"�*�ې���H(5�h�I�*�S��z���џd:�L'"7����@Q=g������nck��D�M: �f�?6ީ�.Z���V�Ǝm�;�ձm[;VǶm�c�c�~�{����e����5W0?�~������5�����;U �$��<&IAq�����nX��s���ކP����^�ᶤ�K7S�&���u�-�(oj�H�Â����Z�q�����J:t�TJW)�TRO!��ZBm�֮�b"wĻUMSOq��9O��z�AYSb�yҫ�����0��G6!���W�0�o>�e�_�0�Q���y��2|ToD����O�l�e�~Yku�J�_���>�� �1��8S%񵂙t�3�Y����B5謚�Ʒ�;�NT�CtVq�0���3�89nS~���78�Ga���v�=&����\�ae��U�����/d*2
J�G;F�h�ٙ�c�ˎ� �U���+�qo��t��ҕ��7�=��w8�\�ud�7s~�����45���+UA��B�JSyN�[VA,+����ދɜ�c����^a@�9C92}�i�R�՘C �dk��,�=��8���c��E����D3��i~Q+M��O?d�z�$A4p��̅A?ݲX���dQ�Ң�����pZ����:�uԠv��ܓ�_��3�Ir+pi/�����wb?�����An���{�=��lw����#�/)�C	���|��8�w<E ��l��w��)S�.��~��t��1����K�jE� �8/X�<�Ƶt���A-��[�-vw�m���Մ������m,ʕDy0˽�O(�/2LX,ui��oc@/����S���L?�D_�_t����~
�S���rb���G4(���&�dZ�V���EK�'�-��4L�r��e?=Y_ǝ����s�vX��`�h4X 59����p�ƍq�(Bj��8`����B�Hq�F	��[�"��CF�i�%Ir�w+�҅är���a��[�J��Qt���)kd��d��V'1����%�	K`
W�/=�����w������7��/Z�0�$�w'�`V4P�vm��Y���LoT	�{�,Ad���"H8$uϮ�������G�hs<Pʘ���j��*���m�j^��]�ט1���-����g(T
��ɓ���-J���_������-���n7��<��� ��#ɭ�S?�D�^g�5��S����@���$�HxFU+�,��C�����~��-Լ�Q�I3�]`�-($P�S,!���ܘ�2y ����9�W��
�.���� �mC��u��L�$��1_�W�21 ;�$5媅�����X&ė)�,K���TF7�WSf`�Y�N�PyS0`�eW��� ��L�F���N����h�t~,��vsB�Z~�a;V����*O����Q���hfP �"*��C}� mԒ<��7�p^��H�(!������l c1e���O�[�U�-�X:NO��X�$I�.=��p^I�����S�i�]*�a�1���ܐ_}���՗�`v]���q���B]+�$@�E�A����kĩAo�?)4�î�M'��5B��]�H'[�*3���ݬ9�)�'�Ӡ`��
�j��}������}v�� jm��+��g�a�}������W�R�A	W,�J�P�g��uJn8g�ޭ�8��!tЗÊ|\~�H|dw��J?T6��L���Lܬ�c�T� ki�[�e��SN����S��3K���X��XO��'�kȅ��G= @�52�cz���)����T���?���ta�Í�tȟ$�SvCC����X�	'�Ž�M����e�o|ܓ"�
79~y�K��T�nj�0��
�^��t���f�%�8��`J&\K�f���o�Z~˄�i�aJ4i�7�n����ۜ��q�ЛM����x'k�|�
�4�?V� �V^�N��8y��k���`��
N��jq)��������o� O�2����Y�]�b�E��:���[Uh��'#�j�#�a����S[`r|�;����r��O�zc�F(���~X�J<��@$]�-�(6��Ƹ����q�¤bh5�T%�<Hæ� ����c���#ل�:�oe@�X_؈$������g�,/��|���j��)|��,�)%��A�W���lm��I`˝4c�<�	bB����<�f�t:;Ӗ���h��hP"v�#D,�W��v�I�7�ͪ��˅��=�@�5���f$F���"�r�x���7�ߤ�	��(�t���}Z� ?a_p�Ո��6ec�v��P5:J
.c��zX}�T�������y���Ya�J�\U �v��4����#*����g������J��{���&�%m#��F�krQс�>�`t�-�V�N�n|'�
��g��2`dKƝ��u,L���s&(d�I֗ϲ�0�%H�J����pS�;�
E���]�{��*7��_���xQ�g����^�̯lL�wN�T�h5L���}8��33m�#t��r�KUw�|���e�cs\��7z�@;Y�n���!\9�Q�������	��Ô�����:{��,m�� ����*�.����,-N��'A߸�=���kGn3g�o�8F����%ޟQ�v{�5��<q�>Ҫ0&[��[)/����e�#W�mg
�ᅹG�2��n �͉�w&NMםl��~$�a�
�Q��4��;�p�����1a�Mi�,����Mk�7�����z�3�����y,��}yeJKZ���mV�C����%�.
����&����d%�mC��4�s��%��V����{4Q��jKB�憧�x�l�5P��ԅ����ǽ�N��y�<��n�|Gޛ�vQB;�^3rh�T�S<��o+�E���2����OӺp������o�Ky\8��O�V��7�|�_�N6�o>��Vp��}�M��yg�mw�nM�s�;"�9���G�E�W�FҍN2#E'W�J�9A��J�}��Vi�)��lj�<��+ͪjH�W�}��-�dfP��P�V�$�Q�w"��r��rv8�M�S7���P�a�b��O��{h��#^��Zy��W)t� ����(.qrQ$�v�|վ���ו�_	���3|�ҵt�b��{;��(�/TҖ���x��}t��˓P��k���&�_�>�%�o9O>f4�:�Q�r�-δ#$%P���Q���M
�?�U?T��W�ѧ���+�y��lsz���T�I?�����j�*��W��D/�j�
n��s��l �H�D��%��菖�W�(�[�����^P�(IL�`�R�����g�r��D��ۡ�/�a��M��3��EO��$�M�h�PE5Jrp�V�R2At��Otd�qd���B��׾���Vj2֠���D�=vĤQ`�@« {s!�1'��TJ6(NL�ґ t-���[�����jN����Xk�����ϔVJ����(TV�lI�	�5֢jdiS�?nK�oҹ��X�R��K~��*�Y��=eQ�a��ʵ����R��i#\�$������i7j���S��lP�M:�H���*7�eD�/��/���%U�@|�����bex�߯�>�wP��Ď�#�@qw���AH���s@���m�.���oa|~�m���V���;��i,E^s��/�E�e�a�۾��3��R}��mñU�p [��H�ݶ��v)���x��3#P����/4���쾏�?T��-�P��TP	�D��"
��mNq<�JO��Y
�Nv����:@�N]�I��J0�hX��怖Fu5���@}"s��p�.\�6�+I�7�:犇�=:��]��b�u�<�X�v |V�Rd0��5�ěZ���}7!����"ߏ�4�)��
"2��6�LήǕy(�%4�է���9 �RT�@� ?�L_����-^w|1�z�p�8M�H�ȼ�&�K{de�Ot�K
%3O�J��L&ws�9f6��Uc�����	d�����d.J,����x0Lx�
n(����$��ʾ������Q��:�Z�HB��Z�{��nƈr�v��ã譎kh1�aae-*� ���@�q�v��G���h�s���hr�|"���6�x^��KI�`���ê	� [�e�o;=@�ILyD�ߪ��Z�̑��̎�jƨ������Rߦ�1$옉���U�����B�w\}wP��,����h��|?��Pg?׊j�/�~��z�_�5c��r4��V�=����������O��O�l3x�{_�{��������J�AF�%M��H����Y(\t���Tv;��#�8?�&'���8\�\K�Q���m�����G�O�_q����u�`GV���Y��f�J$����x�7����Z�P���i�æ�d�:�/����8�v��2T�qy���w�9�
ܕ���,7`�`�H���O�tTI�T#L?������Έ�����G��:�H���THP*���$��p{=��?�̀�b�q��;Xs�$�ly��q�+Ө&ؒ`59�\q<����k?��!V��Ov�|`��c�$,����<�~9�|�����)�U�`MS�%%�셴�s`x�L��������p����0JK���>������pe[�z�k><=�c��kk%�LM,�0F��ƑbO��h+VK�UW�ϲ�a��5�dJ\�Qo}��v}��CZ���N$��Y����+���vxQǽ���� 8^.��ۓc��3��T5�t�~�v#�	��G�W�U��v#�]i�y��!mH+|����FC�j�˲���a��.������Z����VK��6�7�j��>j���_JPt�c~0z.;Ƞ@�޴��,x�I���^/��k���[� 6�F#4��"IȊ��Sg8�^}O�V��D��	�t�*p:͠kt�Sz;?�ħ�\C=�c6rbŞ�C��i4k��r7�LHsꀋ�?�{�$�{#���n�v���$��D�nRR����T��|��DZ�)��u�A��Ҍ��}Ɂ�j������")lVc�(�o�9n�*u�h����B"j��t�����4��<��BP��vZ��/���'����DI��p?ڞ�KDB�>p��W��|B ��Ҫ���U�|u(��]_R��3l��mO��Ft��3��N��6�$
A�hOH�Tقzq��)��a&�/N�����&?�^�}�^E�\�����4ӦMƯ�S��D� �7i[ۢ˵�#�#�cnH2*d�b�P�P����6�4	�SPM���l���� BpL�4UbE���0�q��E������F��t:Y4�T�lHbX�v]�VI�2����R��B7�j�է6)�r�~��«7́����TQ�D,=����͗)�d����ƆT�X��@�(���z��sAjk��H0�z""����e�æ�OE�*^�W�NWm��̫8Sl���ROMǻZ�jkaM0M�^j��ē��7����2�3v�b��;��/G�8���h�ǥdK{����x�#i�����XL;T�6<o购O(�H�1l+���6W�vSn(�`��X�	��)�҉s=��놤X10 +K��:�K�l�Oч��}'ik�,@p5�eb?Jnv���D�*�@����%�<k���<o�r]���0	��!�jJ����8�\56	ꝗ����) aTY��`��x�A��כ����_��']��~M�Q��I�!@�G�9��F:�B�:xO���]PE��R\я�T�Gs=����)�/[�( VY{J�C4��*n#]�$�$AR靗�B����%�f�G$������.{>�́B
�E�hk�/̳K*p;�6v"�MT�!7\D�ʹ�G�<pu���'9�s����#E.�0�?�j�p�cG��}>�`$���e�Θ|x�A�G���Y�"��~u�}w�{�Vu�Sc���G�O1��!�D��L�1<7K�݅�dr''T'���7�R]�5�#Ħ��D�9���G���N�B8 �y
<w	tmoQ����C)���Q�A��d��p��}O��܌�A�������������lT6	����`(���u��x���Ao�͍q���s_��y/�����<�.a{6�۳#���F�����_
wa!�G��:ƪ_,~+�+�#~��~e=1b���-� �͙V6.�i����r�)��'O*{�ة���˱�7�SƟ�Qq��xK��ֿ�E���i�%����V����mZI�ٷǽ=ӈ��r���-`U�!��!l��rG褌l�eCй�~�/�Tֈ{ �,.Ǫ�H��CI)��gO��=u�"�`�%;���ux;]M!��r\:}�?y��}d�_,&���_�E�!��{�'d��|G)<k�g��v �������w%�&�r*�-ZL�F5��	��x�����t��uY~��?�d>�H�i��*v�~-;EU�~S'�~�+8X���0��>4* h��A�v�V�(�U��$�u�!����
̬�ۦ�U������o{޶P�aÎ(�iZ�eE�B�O�[GG�%0S�d!Ts7L��HsV�K�P״���'{���pײ�=O�v�ʡ�L�x:;��97ĸ��V*�±�M�L�{��c��n�]��ve��Dք7�	F�9=���Ayʂ�����Ҷ|���@�֟��<YAD�R�Z$���J1��8z�I�wמ�W;^d��� �R� �l�-�'�Mw?�k2D�"��.I��*S�	�-�� ��W��Ǻ��!���eBF�6otL���9��rm����|�ϰ�T��s�GM�d�vg=��A�h��r�%Xytb9��1�ԯ��31�M��*����mE�X��?��C^��@��g����0;]��]�6�c�tp��������ß,r(�����X#�01]xk/j鷻il,��r�m��  �G5A�~��BA1�y�{dHo"�������}� �ޜT?ܹY�{��vQ`�uo0��ׂ�e��
���`���[
�F�`%��9;Ʋ0�
��{0��-;�b�ƘfΤ�luF���Sj)��?dm{�&���wYs��A����A���BJ�G�1��P-
0�2*����1��&�������C���3������x� ������Ru��
��]3YQ֪,�<�=��*kL�p3Z�v�[ �uR	t,�3J�"�����`,���01����Z��cO��c�(GIs6�S��Ї��U��-�Ɔ�Y<ֶ��li���)�f �UB�A!O*&�d���3#^X��%"�������FɧT�3�W�k����Q.�=��7p�Hr�F�8D�v�J����2���0D#�v�`�n#��eN3+浈:�p'�m
5��Bbqp ��x���,B�h�u!h$R2F�%J��$"�^�_���z�&��J�mPTSR&.@�\�v��y��`k�
�'1�m1E��O�FX�����bQFc�����k�'����@�E�T/$���4��?�e��?V|m�Ѽ�^�H�ڲ|R� �&����&f��0~D|	�G�š�a�!`,���	X�lsz*�`��O����-'�|�q<^bi]=J��]/�ОĴ���hU\�����d�	�����k��yd�N�-���@8�{B�v�}qN�3�^n
N�R�rLu��%p�Y0ֿ癊��'ǘ]pl<9���+sԸ�y��j��l18��h4Ν�qn���p�ϼZ�;\ڀ��|oy�;V���A����i�#�Rf?K'=N�_��x���uq�����?���D��S����������uV�n�V�/����1���T�]�X�|l���W2&?�H,)��8��q�=��Z�R�s�f�N*��7������1�B_�i�X���FG�T�%I�9�O�"��1����
�W����'Bad�:�y�qJ�U��"T�y]�b�f	0��G��CD����Zu'MuQ�4H�ƾ��*F6G�����bV� �7R}���h$�!�V�(q�0�bfR<�"�q�<#���q��㉈rd���>� �̝S.���iѡN�Q-����
�q�߉��D��x"�񜈌u%�E�8�\v�������ڌ[.�Ҙ6��a)~��f �����,$	\����H���s"y+f�����R�fZ}����L��M�A|��xp�氢��eDc(�]m���!+z|*Pm%+a���9?��� �_w*�z(���I=�	}�3��d�����gLD�/F*��p�o����\�Dȏ7���v�� 5� �.\p�D��HO���~������L8��q�iކC��Lc�����|5�[i����dF-��o&q|P�n�9���të6����҈�3+�)̉��1��!�Z�@!�c@�)0]���v�ɥ���W ;��g�3%��j����i�w���݉tȆ���#�z�7_46���=�J�"H�hp�	�D}��3U�ci����n�߃I.�I���q�|��/�~����A �=��Ѹ2$���&��E�v�+2;�d�4+;��v̱	/�i��� g;��Wu �Ur��> ⺠�m=[c; ���(��Y�	�M����`@Hy;� ܓFK-���ʫ�h �Ð��|Y�\.�E�틖���W�C]����$������9���2ۛ�(����#�t��Iꀅ���L���q�����E�!�0K
�
�;�w���ٗRc��P#�@6 ����>BA_��MF�̨�QGmD�T&���Ƙ�LK�0����[��<�i=^$�|=�r��[/�3�+��MD�?���O��jS���Ne�i�&2t�CV�~���|�aW��W��F� �B��n�x�8&���$[�+��p�������KE�4�o������X�<׺k��7Eq�eTnmB�6�6�ʔ�n�b���!Jg�9�#xi��E�Jam����8��H_��D8䑠7�~πN�BP��*��{��Es���:�'O�W3���}����"�&J^��н��iM���KЌ�/���5���i)ǣl!��%�,P���REX�ڥS�� %8_��)������
��}ܨ��*��Xv��!�:<$���!
d���_9(W\�0�&��b`e��u<�3��ve!� ��>�2�������˴yl�3��Z����t`��s�DY����sC"��#���5�N�j��Cy%�0C�� ��u��(�C�!��"c��͙ȗDG�d��_�W��@����P�ΰ,�m���]��yCB�0�"��\B����O��*hf�j��i@�Y.�������3j��i��,�M��ǜ�&�7���'d�+_�7v��(��p���4������E(`��f���@ nPV�h%l�//E��p�O�EN:��q�ry�>f�Y6P
t��S�5���D���th���
3r�,-�Ԝ�:ʓ�Z���9��ט���&(i��,B{)|�E:�U0S
�̙��I�u��6\=�:�vuZǟ
��&D�ٔ��&��dI�<��z]����a`�\��'�
�,,o{�+t��tZ���X�����L��<��M����O�ń1�_1Md���DH�^����&��MT�1<UW�
�L
(�s7�a>��iK���"�
~�;��~��ѥ�%j�
:3rOD�]L)�����9���.�)w�KlJ���Y����k؏���-���I�D�+���s�X�o����4�b��FFn?�/ۡ��kڍ��֓�^�33ۯ'9}�k��h2��z}$.�M헗�[��ZG=Ѻ<B�eA]د�;��(�e�m����>��V����!�c}7��&�����%ܬΛ�>*Ⴣ����pF#�[*��+�컦�XoFYж;SJ�Mt�ә\�Ѣ��5NPľwT[ߧ��6�zs�F�;m�r�vir�)z��;B�bd�@��I�l=C=��.q��d�O�%�rR�ib����	?I��/���K�16f��Q�����KG	��J��.D���(�/6�0�g�ѢZK �?UL}��Ϝ�i��
��C�F��uS���B	Ö�X�7��\D�w��$`DJ��eԼ����:[��?֔�Xm����ڴy$���%�6�=�ۯs1.>����J�bƽ���
s#z�qp��L���K��:zh���Mr�4`��5�p��F徣p~�B&�ư��L���� �)����Q㕣��'��Z���\Ĳ��l@��͇�l��͉*-��㉠v�=b��]i(�F�4�Y�������7:��BXoj�rܜ�"#&��BI�m-ϖ��.W'�^���l�)O4��؀�x�]E�E�{�y���,#����Ѭ'I��]r�&^N$�	���M�3H
:������W�d���<ݠ$��$��8U���J����3�x�9����j5�8�-�@,�q�Ǭ��#�Z�KӇ"wx;̯{X�/�7�\�I���F	�W���3�)oܓ�}AWkY�
���K"�A�FՊ��(�(	�Z�%`�����5�EAx(�-P ��1���̼X��O���o�nΰ��x�����������x�i4bf����4���`�b� �Z_F�1]tϵ�|FM#�_Aަ��ժV�k&9�p|��:��d���-e�%��G�G6|����ſ�)�qAR�P��1Iߦr�bH���ԛ����q��V5�#��$����x�=$Y�"6Q�e��9H#��1�}Z����0����uX�̽ğt8^uy�m��o)�8��Hg��gS`�b@ߘ~t�;�ʵf�����6�c� � G�c�X�|�;�E<�!{+�lj�y� ��QT����"&&
�I��OȜG1�Q3 >�ջfVJ�?i,�@R7�+n�S��DFba�Ux���K�L{�2>�_���PS���|0���9Q�Lû�_�^�L��3G)�/OD3+�e��l��`I��|���I!�1bb[�f�x��G���1�mb�F�鯌�x������p�J��u��G
7UX�iE�D&����@(���=�NR����K���y��~u��'��>��^�ҠG.�����[:k�Ų�6���F=��F�9�"����J$L��2&P�[��y����K�Tu��W���c��}�_G�JTj��N��I!&GR���8K`C���e{&A� ��HM��o��0�;�t��?��iӻwAF��6Vd(x�N�P
1�Mu��������V�)٘."b1�1��,O���o��F���p����["�k?<�vs�iX�A�.���g�i`$�<����ۖFHW�G��L��o���GD&#���ψ���	�Ax\� ��$����$O��5H���K�׼������>#�:QM����'Kv�
S���.5ǥx��� y�J>�e,���(W�h�')�C��A������ͬ܆�a9��x!�获D�yE���s6%�oF��3Fx��<�?�r��L�p}>�;���o�MP����)�I�HCLdo��$P����	�Zjk:�~b����t�&�e�J5 �q�GsITU!�[b�{�R�H��;�Κ���ݎJx�0�ty��� ďN�����b�䵂�inn�}Eh}����#�f$�Z��g���KM>ʩ��c[����̿B ᣌ^ۙ����`!�k_ץ��̒a$��QX�ZN����{	�i��`�����#q��f�*�q����i��0!�nj�)�`|�5~�|�f�s��a�}�ӑ����f�J�/#�-���<4k�������+�۰]P�Ie�FUG��;��G��=.x&W_c�'�"��`$�J�u/�IB"sD���1�";
�0\�Dy��8�=��>���w`�x��2W�0�%��Un(BZ�
ن��J��4~n��@�DK'�A�埱w�{n�F�{{����:P�I��|���4��Ռ���Ԥ�*_)Fu�XcQ�YR陻O�C��D��*��C��mכ"qJC���b�Ϩkz��m�T%wn �B�8�K�-�3�F<�r��,��>��Aw )<��138x�h��Ѭ�nO�� ^��8R�����_��Rq*�.ձ�^�>N�zE@�����b �`w�A�����84,}��ח!�Q�V���Q!g��I�D�BF���f�X�R��M��>�a�I�_KGg�%�<G�&���(A��c���n]0�qțq�t)e̹��h���m:Q��%u���ؙ�/%-�Hr��qͣ��#Y2+��vn���9�����	����>-~*��*���:*v'Ӥ�΋ȕ�Ɍ�EA�P�~90��?1�l�Bb�r�cɿʉe?�aˣ�*=���u�zU愞�Bv9y�[��z#��?����[j�Q����dM`�`APÀ��D:�5=�N�e1i���zWH����`��dZS�rӉ�n���]D�N �̅G㺤�Eļmg�I,�B�&�=~�sD��ع��v��B�l
�ր�˨D�A��C����*�Z��L�z�.X�bl��v�#��S�'�p��8
v��j��od��-���*�����E��[R��~�8�(�}K�q����<6+`����W`iμT%�ZA��kv���nF��1E��@�ہ7�Ēp�,v��gc=RIqF��9(�P��P/���-�IN^ܟ��ӉJ��{���fԃ�ò�ӆ�[�*���4�U��bx���4��Y�G���&.�G���p�C�󎿎�����A0��V����0��a9I�~䠫n��8
8upeF䢕�jі�h�@h9,�R�A-sCm�������13D\x)b?�>��ʐ5�g-��A1���XF%�1[�c� f���5�W��������u�Rh�>{�ƚm�y@���,~ic@������p��[�R����}q�I9� Y7����r׎�ś�Ŷ���V���E��dw�~kc<�NB�������?����+[V�q���ip���n�dH����K�
��m��e�]�)L��k�9�����!��ø�B	�꟩\�j�"+5s�(E��Cb��%2������ᙥ&����~Lr|�fN>x���Q�BA��jȺ-�ܪ�
w�Lf��o�I<���RwI�&@07��ʖ���dG����jQ]�o�o>���[�I�y9
���m=��;���B�\��%/��[{�]���L�����Lnb4���e
SZ�i���T\[� [��rCg�1�+�`O�ط]�n*�ʅRj��IH���Uj@/V���!I;�\h;yF��>�a\wR�QX�[�%��-F�֬���a��]X����p��#{���Yq�?~r;G��c�Y �~K����#碒��eFZ�;���/^�_�8���~Bn:@kV��A�u��S$'�at�wɌ��ڌ���miEC谝B�#�[+ [�
X����_mQ����ɒՔ�ʎ��������t�*� 8J�v���r�.հ(eP����9���㞋֯� �>�,��C�� �ӗ��/D��A9�M��1d:�#!�� �2*�dbJ�qS�>��!,-?��m�R�y���+si��9y�¤d�L�ZǙ��n����A��Zeߟ����M6 f)�F�+{��a�s���6�����T��=!ݲ�a�E��6��� !�y:rJdoN9"�9{�1���x;m������)dMR"�Ī�@슲B��I*���J�f��o�b��f�j�(B�]f�U��t�]��e�C^U�ۖ��I�U��.����Qb������u >҅D%���ff����7ճݖ>�^�Jg�`ʀ�L`DM�����z: �5D�:�io"�i7O��Ca�ו�c^���?�d7
�w6��K��
2c,�$KB/B,ɛ�ys�4꿊a�&�N��賦;r~N��j^�Cg��䌛p5��q��߿���s��d�0���`��a��ެ�c
fDy���NA{̈́�\%��"���T$<P�瘳cQ�=��4�@��AѰJ��T�V�S��Z���B\q��}��`���>\�&o�D�����{8S��qlƁ�Ô��&�I�ᡲ���F�_B�cؠQ�l�W��)���G�]�2.�D˞@�A{��*c�q o�
ֈx^|�N�3DUN��	(��fR9�g*h�\C~jT��|T��VE�n����\w:����,*�`����Q��Z�1**���a���D��F��b���T`�HA���JVY������U�Ib�
\a�G)�jG%ވ�#غ񝷻�,' mF���p+�^F�JX";�Bih�Q;mtDv���{GA�e� QQQ'�}&��OK��/��>�SOǳ,9KU&N��gp���@*� ��r�Vq������]YqsTõ��ez�1p��'Q�g������ 4	 t-�j��P:V��s�+����,���eXf>�$&���BJ�T�i0u�P�N,F�=�-lg�\&8��T�"Ͽª�;��{(Pt^LX�"�']��p�E�������-�����R�O�&����Z��f��(rQ��CU0>'�oB�,�eϗ˘E�Kē5*�u^O�z>��*���Ka�x�&����kP�Rv�6Y�b�RI�YngC
��HW�2f���U����|����R�	�U��EN�m(�<]��q�7xl��̝r��U��|��v��m�I��ajdR-�p�.�Ȣ)��pk�T���S�Qġ��Ɏ+�j8D�����5t�8�Ǭ��Z�S'��F��<Vy��	H�%��%�f@l�m��S��3h����+��aC��K.�<����G�|���k�S{dj;b�!
+��#�[�Vp��4�[Jʣ�@���+.���}���"��+4�冠5Zh��q�ʨ���3��GQ*��R��G�B�<�_D�P�0���-���jFA�޶g2-f���dw�s_�W�[:���4�T@KL�]�&�{���$5�'�|��Pe���&��$�I;r#���X-�>�@��Ɛ ju�?^h?�.���Aݎ���Dŝ��#�IO�Y޻{'�*d��c)$�^_w�?\��+!�*<Ȫ�ɸ�(ڝ>9���k㖛ۼ�H{Ag�R�t�T�����#+��H����J�1��f�7Q���ضӐ�ő�M�o�E-(_������|��ܜ�}�x��\���G���?,��(�HQ���*��h'�Rŷ\�`�����bɬ����ԥ	lj�:2�lx��e���������7�uM ��7OXH�|�FF �KS�ߪ��y`�/t��&P!�f�F_ָ����]*�&����K�3�&4�'8�̍ل:��v]�������/�\�z�U1̙Yv���&�~O�
7~!�8�9��6Re.�)�r((Ħ�L��LM���F���r���NM/sl���(ML*��c���)����	a��ٞ�?�-�y$3p���H<Y?YU�ʡ��;(���\���4�^�.�F�YU��=1�Kk
��?��ψt<�𐤄��M��Ԫ-0R�GaPq��<�[��,�p3��m���!G5������P��wL���~�V�S��I$~*X�r�t�k1F�U_R�����F�/��6(�����'ђ�E@e�uY��K�ӌ����5ߖ�[�z/:}�y���rm� M7�L�QJx���o
�I�ge����ֿ���"��i�LP�\�gx^ۊ/��l�螝jc�[�oJ��P�
�I-j�V���F���/4�y�\J���s]_�@�ǎM�)��K?XL�Cn����@L�%�l�4hCarh*�~'�b���N��'�$�2�\.�cMʒu�ͻ�_��k���0����z�%���̬s���g������J��[�8��D�&en���S���x�M�N��#[������n)r�L���Vֲ�<|T�;S�!ޣ�4��)��S`�f���>��1�b��Q]�!]N~�����,�^�YQ�T-�8M��ʛ�2�\�N�딍���n`򏏅sᯣ�*�v�hqdN����t��)�Y��i�uB��=Ǹ���8��Δ�΋'<?]dͨ�b���ݭbsyY1���l�Ѷ^�F-W'x����S�1'�X�I�~g�FS���-0�#�Hee�Bz�Q������r����C����I_3|n���S�T+�S O�F��v�m�������4��⣔�Q(9�Q�N
�ܢl�\s䦴{'�~V�����4a�.ʲm۶m�˺ʶm۶mu�v�mۜ�yg���X��+���k�����N�X��Q'S[�I4�c����jK�Ӭ�s��X͊W��hHA�H��)$����U]�@�>n ����H7�gQ.�4r�0��|�,ER�g ^|ckm�J�nЙ1�X/#���ry�q�|_��*�@OrrѤ٧u�J
%��D�R��띑qo�־�;��p�i$Ⱦ�v��K��&J�Q��>�#�v"��f)��QJ'�0}$�
&n3,���o�\�|φ��,������k�9���@=A��JA%H�i��Y�05�`<��j{4�m��_���W.�j��4�)V���=@Xn&�VI�H�����w]�t���D��X:�|���v���m�I3ֈ�s�?�U�z?`�0�@�[J������KO��c�I2L�)C����2����
�)S�������m������5���D/���&�����ad�R�Tr��QM1�����m�!��Q����iT|�Y'#>�����S�I4)O���WF��Y&Y=����4$v!u���<'�ɪx�J�����X�x7�����r���58}%��L�4�cIL��A*�J��#���G����!W+%4�.�AK�'�;���Lv�Xxˏ���7�K�W����'��: ��sXqI�Ѩ\QZ.I�F�C��S�g:��G�-��B���=p�pL��s*�H�����=��l�io��B��o�0`�GM�0|�2�~��F��)��ٔ�=��jx3X��]�E���8l��U��#�Xf�_�Gӄ2�S
CBa��T&d"���Ȫ�hF��\���c����v�43J�S�ڵIn�xe��>K`H��`��� ��M��'��T9B���c1lXsG�f��0�u]�;{
�Uv5{B���A�]��imN�Ji���L�}	�Hk�ě��6�-��  �eTa
� ������禙�4�F���VDo�!7�H%i���@�kҫ±��;�0Z����Gf���-���3BH�'5�������R�R�@< x�z�Z>�.���\$�8mz/4^_����v�ȃt�����q8����p��s�&��?^�d݄6��-������Ǣ8�q�G���|�Ā��=���R�k�om�v�"*�q���>|�ds�]�m�M�C)��9��&4J׌/�;䘀 �������@�2ͪ�'��C��n�����-�u%��+)e��;���5�]��;�6�Q�}��R�D�v�ۙjxxJ6����Iv�t��2I��bn�/�@�4�۹������伏���[�������o\�!��J	�w���x~#O�Pw��6]�[�k1�g����F[�v���"I-�Փ ������
R���G۪ɸ�͇�KiOf�O(�`I��Q�P����=J�a�G頇�����g^� �}x��W�������p*���w?��:�Wœ:X7,�mA<��|3����p�fĖ@�N��h���o��Dw�xQ��hԺ�|$g�S8.D��%7XB���HƔ�\X�~�}�L�&������>��k�p�Ҁ���Qg��5�����)VN��شઌv�ܐ-��uCo�8�=��w:�>)PW�ؔ��Շ�LI=~�O��J�4J�{v�����@r�\)��H�������Ժ���L�f�3��f.aH�x���G�����P�6�ma<9$�b�Z�2��4�c��b�Ҍ΋���9�j}�q%%�8bR7��54�u������g��'��|@0�����:��v�n�0�]�c��@��/��ty۲H3T
#��RX�ܮ
�@�;m�N]���Z���N~E����
ձ�7Qi\P�8U��0A%���Ѐ�p���&���󀱅E�e��C>op��v|=��2���_�QBr�?�i�n�;���ND��GQKE.��ⲫI����Pe����賮;z@\� ����h,�A��) )Ƨ�߻��q���Dkf˘27�����/��=�1w;d^χ[�����r+�9rsJEIS5�D[�w5|��^����#s��V���*bmKH]�A`�9@e����׫.̀}���q]�����m��̖�i�mf2�-`G%�'�\u�p����������N���遯���'$��ɡ�k�?gDg�\K��z��M�2����xo�έ���_���!�C�P�r���kH�����VnШV[�1h:���d���́�`#�\2u� ��ƃ�r~یj��<��<�0X���Ho�|r�1=$�iS!@���X=������/��d�v���
��L�����D\���N����2�z	�?��a�)I�J�5�m�h��8�0Q�(#�AtT��MvT�i����c��%ŋ!���nX[ikݸz}����|��7 "_�����7����2?�DS�VK�=-��^[�++s�1W��I��m��V�7^�yp��)��5�Q�}>;�s�]+��(Y\�K��ȷ[����p���LM|��F�6��x˛/ۯJ_y�����#�9�d/Gf#�r�d�� �0�1x\"�l�(-(����1E}�c䘹�zn8���\Q	m�<x�&wk�������v4:)�a�a33��&\o�8B�<a��P�oo����]��9(��2刜��M�1Ll�/�%M8���ؓ��WD�pX�[ri���*�����Ǹ�����Q�Ո_ql�+�i,4�@�I+����IVycp�z@_����!�n��9Q$�d��R�lK�ؑ�Fk���&C!:�O�*�'s"�x�8Mmyh*��X 6(�|���[���4�a�����"� -��1��1������(t&)��j�\�Ѽ���W�KW�o��Ffr����8��a��#�u<̖��Wt�xΞ�a��M��>�� }h�u�b�b���&��S'�,y���O)�(�o�v��{|R�x�f��A��4�d��{jx���>��u�k�$,ɵQ�ou��v�-r�3����ő>aQ���jS�5I�S���ȡ|��&�d�7�Re,�A;�HŽ=�H�c��e ��i@ҽ1�|d�^j���x�k? fMԲOf�dln�m�#���:>%C}��2��]�Aw�
�k2�g�[�8oH�	5�ݔms����uc��.m�������4}LU~�ZP�+��+J��F�A����f�Q���O���/�Й��c�A�u_���k:VF3ڿ4�?R<)����rd�gV ��*�x����6KtZE^��^P�����Lj�d�j��K�՟CȆ��;�?(�S�M
��&�̨V���p���]��'��J��M&�JK�bQk��X�N�F4�m�o�1>�:}�_O��k}X��4��*.�i�)脣ȿm�\ANm�䡄jK��68�&>b(�l�!��N3#���2�řIB<�b�����Yy�l1
[�:D�`k��b��'��Pn���Ąq��&��N�d�E�YKsS�B�?%Y9X?���-�닕1!�?*Ѷ�tY�i��H�]���u��l� �_�e!/\1T�ˮ O���]�uxv�߷�!�8�'����ʵ졡	!GT��Ү�z�t�%�a���C�T�?�45X �=X֡�
]{�v&9�Z��������[.�ϫ&4��5���"���r)xpv.�a���7�h�;.�'�am�a"������V*�.`t]�F^F*	���T/OF>�T|��Iad�.U���(�GN����y]�X30�MX��P�7�\zQ)�tjb�����#b����7g���Ҏ���Ɨw�:,�vvڻ��8y�oQ�A>�h����CގG\A�Js��)�d�>���Y�fH7=��������RS����|�Jw�9��<������2�g�PN�~�ԟ���|��B��ʹ'lz�&0x�~������ 1OHO�HA�h�rt�o9$�'��r)6�X��n��s���^��%I��&�]���7s���b|K`�p�L��ŋ���\�vϪX�y2E��ڌ�C���?�]��zL2������#Т�K��Et�N�j�F�jMs�^�+�x�|a�mT�rD�4
;T;~.��9� �f?q޷����v�&ʒ9�M�&��h����#�i#��6,����;ֲm��)�M��<Q�������=��6~��FoF�K���=O�Y�������-X-+Q���	<��<-y�mK�d��� ���@�:����?D������^r-��g�(
�g�	�M�̌ڝt�Μ6�˟]�.���y5�؛���� $������u_��N^�돃�B0!���7(�L��8��nė&\gF��vM�������#��f���T@
��b��5�p�᭗m{9���j#�<��m�)�Dq"b���@�䖜�*N7,�9�_����R:�dyDq��x���B�gBK|��/7�3��@�p%�r4Xd��	��|��&���
"�cw���;ݡf�(�\�<�|�r����Ʉi%7�;�0��Jj���G&6[�bu�`U���Okd\�G��K7�.�Y7�w]u����1�=��#Sa������C5TQ�̑*��Y|��v�[��|?��Ķ:� �*���T�`s}�����^&�H���B+�'\��� '��#b��eT�W���31ZՊj�oA� �߻U��" �����b��;��
��ق�J1��y+��k��HV^�D�`�OO+g����Iz:g!tj�Sw���k�.X��zH�CN5��M��i�æh񁘂(v��Y���p\���"�:>;^��%m��y�L��SI�:��ʂM;༬Ab�(�__�L^��n$�����f���F���(N�c;��j�����D��3���l��n�=��^�/�gG�c�՘�3&�~��Ҁ`����������>F)���1����H�y��,q�7�|j�� w	';ʟē[�/�j��ވI�f�;KW �cͤ��I�RZ
��#@�7�n"��~X�Og�T���5���sXyf<����=�I�6���r�rK!I��izt���n ��=/a�^*���5� !�X�r�@A�?�X���1u4]C楬Q�+�<9W�����
����<�9T@�x�bs_�V��n[�*JaU����1U�m�0y�o]iKA%~��^1���^�����鬇�l~'�p����at��o� L!�<R�_���X.��Y]z����=�����ϗ������O����WI���O.�Ĕ�t��9�'*���۴��v�<W�ckM��1D/;�r�T��{ӏ���7�pL��^�� �
�G��D�ϩ��vʻZ��7�X��%�j��Q)\�����gy�[ʾ�-O������$1Y��Dg<��1q8
Y�ԉ��JDl�2h�$yώ��h��U���e��5�o�C�>�|x=Ke�ъ������ܒHI U�.��u,*� z�r`�(x �`m4`��J��Ӏ��1�#�=| D�^PuXW�/w_���&�?o��L/�6im�>Z���,�ϩ^D8�*���_���b� R�(���>�OŻ��/b���6P�V
ȓ���x�樼����n ����u��I�Aʸ�r��qi�@Z �68�g3�@�X/� 1���!E��À]�$uxyi��\���b�<I�5%���  �1չV��u +�ir#)�����+ؔ{{�i���.�ʊb	��ȸ]��G`6[Y��y/q���-x#��.t	�!P��m�2�Ur"2������=p�?�Η���&\˨�����1Z�j����(��%��-V�'͘yzѽx n�MH���ج�����i�KX�u{���%��tpDz8av�̍�x��~_��m5�m=�v�����W����HI5�{����>���7z� �mV��fUcԥ���S��+�@� pF��;����sY���p�~�����͉v�Ѱ?E5X
V�86OE:�j��q��>�
|�^x�Xl�J�b�eAo��~�w䖉˾q�z��+9*Ϙ�̉4�e[A29�.y"�I�3�����Z�x�\4b�G�|
@��h�E ��
m�V��F]���G�(���~��M�y�ܠ���]�ɟ>'y�[N4b\tԞYt�o6���X�c�qs}�'-���Uf�}��N�ed��W�x#�+�A�3��������D��im�8W��.A���]\�H�/%1z�e��!5�gg2<[^�� �uZ�k�Rp���� { ʜI?��'�:#Q�Ct�(� �$f�Y�f&���y�Kl:Oi�ب���*t�?��!��+UWdс�m߽W���N��6�BZ���w1l��2�瞃=]72X�G�au����(��^7OOJeӃ�-��Lx�J1��e�7�`c����'ϟC��\���g暎�;6��q����=��N��:XS��Aˆ����%$m%�E�`i�I���A;;�|�t��V�o���*�@-6�fb�Gb�ף��7:��:nZ�}v��Kaeɢ�.�8�fj3E3�w�B#lr�v�,t�-��o�P�e���u��9�s�i��H����e�3�5DtkP������W�Ϗ�d:�Trh����%���J{ZW0����U�WRd���e۪+�����9'�y�=;��!��k�@J'�|^��vm��������mX|�r���P�ј��Uaֶ��@���`��#ȍ�A��#��mJ���u �o!:\&��K�A�i��!�3��"b�~��B��^�ol�;q/�� `��xc^6.������?�D%����^[�f�.:h����P�M�K�MpAK���7�����ȴ6��@�I��*x-����U�~{Z�t�%$#$�A�J�,��hϢz~�������V�������*D����}\�	��BN�L[{��oV��'Jg��
+���3��r�;����s���HFG�_�Ǿ_(���d�"�E>K:Tɠ؀;;|[P�;We��#��%|N����[�K�����B��F�>��6$2�Vo�psV��"�����(Tʶ�nN�]��[����]�!�`Q *�R��B���Z҉�e�� #��xt�� �C��ӈV�.�	��n��̀S�B"��y'������>g��ȱ�A#������y��gO�RN����4{��r$�x8,L��<��G�C���S�r��wp�Ak���>���U�g�X������u��9k����
�v�g��]Do�2�� nP~�!3�Z�����6z�f���c���nCh���跧���>�.���CYL�I����v�n���<��%��Ҹ b�TmtzJ!�[&;����m(��SBHI�#������Od��ٲ ���w��V�mh/�e��cF���Wn��,�ЅKaƉZSL�
����&��:�PLKO�ٻ��s}�
S}=�@>Ok��������=�N���8�9  �^���G���XxX��1��K�Pa��bJC�=���@��ꔂ�� �9�F�T�_n<�����Ҵ�a�:�=��k:<K�y��ލ�p=՜��ax�*x�	��{��h��NN(���#޻�ݗ���.������HU�4�O�,y��Zf(Xo�&�Zt�o���M�b��x�B>J����4�Hx����FeP�+5�:δ�=�~�G�<���b̿l�x-���;$ʟ-R�\�1l?��KDċ�}� O�������������%3�$�[���w�AL�����Zݟ*g�XSJ/A�4Һ�HB��,V���^��j��6�NE>C2���T�d(��/��l����e;ΈS~G+�����y�a�ݘ�+pN�p9iAj]�ޘ'B��H����S����S/b&8��bh>?��n�A�S�-�������o'xk���O����R�=��Y��급bE��V��"	t(K��QA��Z��Oz{�NX�"p=�D߿eɟ�낈�l�?fT��B�.*�)9�>��@	f~+S�D؍ ���g*�:	Ԧ�X��(K����}�N�L,��(�҉�t�y'${X�q#�|QG�T1�
Ts�Hr�G�����w��wg�.68��s�0�`�8�gU4��t*5��I��}��Ҏ�w�v;�त�!ss
�C�q~��ٞ|W���3z�ƎF�Ţ�t&��Լ��y��=���g.�>yA^C���F����a��*r�e�D&ḘR_t�ܣ��da�
�B��#O�!@�:F����Ho㘋 ,�l ��Qu� 5:��q�z
CCC��&�>�i��X��TՇ�D�X8�hJɳ'��3KsQ�*�,�؊���C,��h�W��h����z?��
��=�d�?��tOmx W�ad�Ζy:�9,�u�?��ť$Qч���~�(������"�Tp9��	�'�f����F�����-�m��M(p]%5��6�Pځ��ܷ���Q��k�-ؤ�s���B4�ӭ�=���ciu�b0lc7jS�wBY���{ o���xN�(�ϸu&�����߼�����6�����9�ޔ~1L�����v�2
&����rή�,����%ri�L׿�n@��Gq,8�Y�aOO#��uI�A`g	P֏p�4��E`�mq�6�-o��z�s�f��S6\R`CK��%&��B�f�)N��tUAe���K�Џ��Y�Q	�َ5{R=x�,KW(=�1�^���M!���Z��e���O����������S~�Q�Ι���&�h:~�c�P��e��ħ�ldԮ ��X�{��9�R0e�r�Dg�?_�����j	ȳp�y"��$M$�.��*d�S�x5��!lL/5�H�vLD�@�US��Hr�@�8��5�Q9]�)L�H����b�jA�|Z��af8"TUIAl).p�r$!Ȳ� ��Qba���#N,~�����F�������G%цJT]�=I6�= zSհ�#��Z�K"�x�O�!�D���TR����|OS��C��+9�BM��VE<yhg*��Y�w�7�u9`@B��,G⭬[���4�2L-�w%�Vu�J��N��U!�}����Ĉ.��ĕ�� ��&_v���CO�������M���Y~3RU���J�F&�a�� ��d\CM��?��U���܉�֋'�ʹN��Cim5;;9�z���Fî ��Z�q�;�c؇�&~�#kI��X�A��_����q��fK�(+2�W.="�Bc9>|00[��$�v�q&;G�E!9[�f���&�{�z�+ �ciA`����!�LAX�7m��N_��{]�����X䟦�DuǓ52\�_�Il����Q�,||�1�e.z@�AE���������!c'��b��1�fN֣�<j+��F����ȸ�òDdi'܄pj��-4��<�>�������_�M�8$b+����A�Qx��M�:Z����6�a�����:\��#���%��ώ���I����9�M��K��A@p���U�i�J�:T*]F�\Jg0�P�gp �������5��1C�ּ-�l��r���ӶoS��\��O5��4b��&�ĸH�2}A0��Xh)�N��g���1L�L��θ6��0e��'��f���q��bGr��D��1��q|��| 
G�oZ��dkhn���#a��:\O{�w+�n�:�"��	$J1F�Mіl�X��#oCCs�/��0�z"m�Bۮ���E/����g�]`Q�_/���I�@��wIn�ߣ1ǯw����V��Deep-;�<�'p�S
��m�
�CJ�o0�}�w�Z!c*|0T�q�t��6�n������Ą�
<��0�o��@��vG1����m£��MZ�tŘ�VYg�����NP��4a�����o,(�|�l?�扡U�l�̒4�Agq�mL�)��XN(5vF�~���H��,��D[�*��.Kkn��%��NޣbWKU��+0E	"��2�nɵ ���U��eA�wP��H�τa��*qZeAI�o�y-Z�J��S�x6�w�l�G)�7wT��d���G�@�K���0�� �H�$���[ƙ���I���.Z�TRЯ��W���d6�(�8x�
4��y�E��Uta58~u�0�e�-�#5t�W�NBw�����"f&�8��If�n�[���
aǧ^*4��@=�jI��BH.�K�I�w��6�� Q���>��i�2�cv|'L����O}��O�k��m���#�X�`
7P]-E)ܰ+�ﯔ�oR�#�;ht��ۋ�@!{����O�U��gT�����{��� ��l����O�s�����bq���O�?�h�~�������/�=�����y���2#uY��P����G�o�N5l����#���<c�Hvg]���(A�Xa�M�\��n� �/�+@NՅͥK�Vx~�Wq��/�������lnF'���N��:h=I���M��#Ѧ�d�$V�}�G�t|�9�OV'1���)4�2[}dr����Sw���L��D����>�d�Ң��9'��(��J�~, C<�A$�?;Wǈ<i���Ґm!���l�!2O(JHbK��[��BGȌ�Ӹ���� ��u������,�ItUEL3�	7�
Vu��/�t�uxfdNf4D�"A�̊���p(�� ��rMZ�`5����)�'�5Mc�*z���m���ź�f�F�`���L����L��'�ݎVbt62�`%�0�R�[8Es<�ۘ���4D:�2�M Z.��
�Y=��rf����ы�� � ��1�["�Z���h�|�}��؉P�b�49KG�����-o:��!�����͔�dD�qj9s�`pn���A"7��D�m6�acy�䌲��G-���6���Ff�(��_����v�/�_�H"�X��$xP���z\�M�D����L���$�^HE~��p�����Б�(вO�Ц�7E�MR�Ӡ;1���rp@�q���ܧ�n�P�_�\ϙ�O��������K��@�q{�o���.�`�ޞ�@��\���n.�uʉ�H��=�����3�Ӓ���� �F�!�.	p�P�h|f���C��\绨m[�e}�3B�Á�KEU*�.*��22(�w(�������A_W;'��F�a��е6�_0��)^�(8o-8{�Q���U
&�e±bR�}a�fJ�ɒ��������� ���t|Ц<]�P�Yh=�I�w�ͩ2�m)��$�z�'|Di�̃;Hj6�����b��IWM��h,��t���M��L���G�'c <i[d�^�g iA�S:.ބR+'�d�ͨkCH	ub-�ȞEUWqh�`�B�޸�#ح8j?�x�_�C֮9�s��l������yi7����(eYbZnYi��2�(W���gs�: {�`C�L��-�Y'�4���b8Tb�ꢷz��Qkb�x���o.*rS!��v��KaVK*n��F�EKrx��×��w���/���_��{�U]�%E����̲���vdZ�U�1PTD�d�i��&�\*�<I��A	�L��j�WO���V��i��w�������I�g񈇉���h�1ˤ��O:��F�V�f�������F�
Ak`{_��`]���cI <?�_�^����,�^���/`�<>�t3+x��݌�I16�:m6���:˴P_fF�q����6Ayb|5biְ�9a�Z�=�Ax�������!mKA��+m�����g�}^���`��$ȤgUVFtKY�#Y��𿲰j�\�Ħ��8�����;L(9΀Gc�6�K�nK����%1T`j&�w)�6�����c58l�ﶈٸ>�i=+����5�A���&$>�`]):��h�T�E��m��/�b`B���hch*ͨ�w ��Z
:hIs2��Ѷ����/��ѷ���١��{�
/m�t�����^2�@���7��r�iu=�#��L��/�`Y��R���� A���4���L����H�*񨙒��vC�t!Ғ�f�*�HC�V���[�i�D:Ӭ�3�����	џ��T��?�
��2�߰��]>�{|���h�R��W�(r���[ј�$���d��/UP��⹲�����qcH�$/�1��G=!9�V�9w��͈QO*��0�F�)��XC�������
���Ž���+vz�jx��/��q�'����b��
��s�V�ĕě�Q�1?��JEDA�/O�A��H�K����l���Յ��\�`QB�/T9~�9W��Z��!O�~�UkX���C�)]b�tG���e�x�055b.M�
�˚3�{FT$~]"��,XuI2E�E��]���?&vU��E�N��zc��`���ø�5�Kb �y�|�/��h�7�ɩD:�H!h��H��
�`9z��ҽ����y�<w��6�ߴ���x;���m���QDMjZ�F3�E	]c�Y�qa���]�+5�9�g�ѱ/.�`o��)��p�����"� �g�l�
���=�h%,����Jbl�mC��C����b%YeR�!8������i�7���T6j���'�:���c&
�=�����-����\	J�g��u�l�1�X"�h���ɨ�P������}��o��S�S������O��ӽ�-��Γ�|�7ѯ���ʩ�������qH/�lcl�B�R�2]I��s���/Cc��WAj��eK���\�|!��R5.����+�°\~'��H�%_S� �l%�A�3Q51$p��6�b�<��fW4W���I\6�<�luO�����z��f�T��r��rxh'2O���M�6�_�\�Rb���*�?���X"��K�u��a�&�]�ɂ���dqZ\��p1�E΅�]8DU}�W����F;\�P���Z&o�3b~�a���tt�,��f�n��o��/A9o0rn���NE��q)�QQ���q��_�t�%�Hf�[Z@`�ʌ�*��C-'����s1��30���T�)�f�>�h7�$	#E�Kͫ��S�~��c��ib�-����Ju��!
NJNR���\�4T)�r:x�A%^ ｦJ�'���Q�*����U��	C
{Zx�N�\^>_�עUWN>���d���_uR�ص�ʬ����S �U�e�,;����]�Z���	�:�G(ym8�3�"t\��Â$���Ckz�ڰ���N�Fb��&�Q�Dc|�#�B�n��9������~��n�Z���/����P��Glz�@���W���Ӧ�V�V,v�u�~�o�|��R�ث�dF��T�r�J����SF7V�$��x��L"_|���]RLJE���'��/�Ə������;]F8����u`<�ҿ%Ko�k͋V��jË[��_��Gm%�ltVUF��m���l�Pu��ꂌ��8%�2fU{��vS=�x����O�ŏ�~����J�/쭯^f�g$k-ju9-n����]]�����Ĺ���&�\0�w����OnGd
�U%�\$p�RydXLg�V��qt&�cY(�޲�~�95b�b�Rs`J�U���|��Ej��%�?�j��Lr��������G�j��ߕ��U<����y?��6ޛ�3p\N�~�Π����"��N K�!�ē`��6Ӡ�f��%c߂.2���0�C�ڑ�4(E�K齶1����0�ึ���3�Y�d���(���e�B��ȗ�Z����tF�P@�4b��"iq	��^yX��Z*3�D���[˘*��0�x6Ϙ+u2���88��"ܕ1yDlڮD�	T��2�qH���hԏ�.�����v�'�6�����Դ�k������q�w䚱q�����/��@z_��±�&��2���y_���i��C�`l/����.g��u��m��ۂˍ���_�Ȣ�g�?J���~M����~pBLɑc  &Y�55��4[`a=�2�d%���K����H��e����Z��<���i5<��������6e�C��źh[%���^�(�.0ľ�/8>�y���:,XSEI(���"f*��Cmt���op�E�m�tIdx2�tf���iK������r�8�P����;$��m�>Jm�0aȰ����W�N�������gb�o$���^e��G|���_����(}�c��h
������'rۯP���gG^��V���Kh��ː0uA��I�`��w'�0Γ�I�NH�!t�"L�!�q�^�UB^=�������R0 �:u^Bp�A��� �T|��B��_6���"�]F|F<���C����cv��1�Uwn�SK���
L!��QFe�w��Z��d-W��w J��y`��5�g��/�{N7&���;ǇjF�~MW�ߨ�EG^�E�	=5��V�u�b	[k�h�IM���� q�b���i�f��o�J�ذ\�r�ɤt�_����j����Q��)���[��'�J9�/t�M�5�u��֚�5�xN#ڇN���LF-<z��)����9lE�v�!R��� T����קBm�A�u��A��+g3I��H�d˶�$F�G4TshmyE���U���Xa�Ji^7�$��u���t`�Sj��@��3�Ds�+�G:g��O-�ǋKw,�L<G]��@{��t�}Ա^tJ������5֘��3]�%��7Re$B�!��nH�e(d�RQ�~M��Қs�)�F�%�ϩ�t����|\��Zv̻O9���a�_��GE��7��V#��U+�Y�S#��І���"g� ����H���b9ޣ�T��B��w���^p�k�M�KcZ�J�4Fl��&���ʜ�T�Ra���],����h�ϘE���L����,���r�O;j"w�ę�#�t`e�9��p�(���%�ɷ�MW�F4�S�����f�d�} ��)?�o�q����a���ȧ�f�Q�Wz�lͫ����a>�m����(Ċ��U�������[�:a�E\�^F����:&ǌ\�d�X�f� /���[ڙ�1��l|���8�&��e���U�>2h�<2?h�s����:W�k�2��+bdP@�$�z���m+�!���� ��
)�{���kz V6˲�����HJ1}������崖;�?)�HZYLX\y 
����
#Q;��w
�Ȥ�Đ������P�>�����04��(�o�f�S/?��]�>>��I�VG��B.����TO
��cܻ��r^'^�4lm6����pyu`BIv���C�u]^���O��x!�]�<����A�ԆQ	Cq�~C�a�ۮ�E+SN��l��ʧ�X|1P���/U"2-#'��(�\�q��U��R��Yu�p;I �^2���}��@�҄�y��s7���`�B
O�+Y��	}qJQ�*�~��ș;�	?!XT�%��d�F584��.-��+��&1чi:���}�x�b�0����b`���_[>��\W	=�Rxsd�C�C�����y�F(I̠�z�fX��d/��H\�[��0nx����w)���Z��Te�T�3�!TJ��L�]ؒx](�~'lM�]!F�7}]�;��3�ى��M�X� ��������ń_D�E?ulv4{-���,+�P�Dk�I�qѳ%�����IWQL7:#��q�H����VCn�4˔)3��Q�d;�T�H��4�qs�	\�p�#d�i�	���kԔ�RV�49����xx�:����҆�)ep�ԬV�A��옣�VD���$=91Դ�T���I���#Yw������J*JB��2�8�Fy�D�oR8���x���Y�Q5�Ɓ�D���޵\U�#b�Ý�0X�e��S��}���~�1�f��]���:cZ[
í׏�Ж�n��������=�8������(o^k���;*Wn���)�6�!F�ɺFߒ���ȫD1aSX��f��B��e����v�D^�q���p&�oR���[.��zO,�Q�}�|]t�D^��d� Q|���A��ș��j�"J+@K��c�/�D�}}FA�
[�b��� jg˼��{�K�)t3_BQ:,�*W�b#BYP�y �9�:�����=c���v(X�gU��vwT~)�#��٘˗�Ƚb����o���Ǉ�u�a"�s��I�MH� ��(�gG�����r�|=D��!����m��/����k]�M�f<�`��u]-k���+��]@�����s��5YN�/�MӇ�@���a���[6���ضe=�wO\��,��t�w�ት[p�]����b�v�e� ,x����BQ�c��s��2�2��֣Y��4��׀B��f+��END��:U�� ����ގ�w_��Cc�,�J�at4���$ڒȴǹ-��7˥&U�Lo+w�8�X�gS�G8Z��S����[aݥ��Ҙ��lV��6��4��>.�̹�hO"��@�"�TL�+(��`
����l���ݎ�	�Q�G�c\��O:�S^��Ov��9��+wW�;ҿ<�-��
�+�o�q���Ů[�o��3O�ۏ:��X<؏���<�۶��f��8�7�Hf��t��=�K.�]��Q6e2�i�N��	��w�qii^��bbtm�l��E����U��w��=|���qު�� ���td[����ɉ�.aX^8��M6rME即3h"p���u�=V� M4R�=���1U������ʅ)�xܛp��óhO�p͍��Wzz�uҀH2U�]��3������/�|-V���R�:	� n��������Q��a�@{T�H��������gᤣWb&�C,Ӊ���I\��`�:��2f��it�%q�G>���e_TKw�1l�2�n�Fru�$��t����o�[ଖ���8��=q�e���y��g�n�b�jካo�cy��v֮]�E��cێ<~��O��v"�+���sq߷��1G�<�'|��/�T*BK�a"_�]�����@(pZ�i��%�d�Q�i�1������W�5�^qU�H�`Q��	ZɃM� ����dG��0�:�����G��N=��?���Lg7=�h�5����8�w�'?~��:4%U����t�<Z�L��D��dkg�^+@� :�')��R�(�H&T�����|���}��3��:׬y�;�`�=WrL�*�&���+��?�W\s'��b�R�l�Ma2�k.�x��9�數���߬�C3wi�"+𱋿z��m��F�h�_��T��8`�(f0:2��c��a��
ֻ��r+eh��@�>�
���T� �5	-)�e����Cџ�J��C��2�w�XCCB�|���yK0�c���H��ʐ��F3S	��������cr��SJVCf����U�u�-���FK�M������N�%b��.N�t�G�8��.� ����!�+bէ/���X�A����YFcf
�����Btu��u��+xf�v�z�]غ�������vQXuizh��%�i�1�7���v9D��H��§W_��"2�=��rp��=�p���4v�ԫ���P,��?p�}�Ԥ����J	r\f�-� pv��#7����\�
�,�grH$;��S���{����X�d����88���ߟ\�l[tC���N�SX�x������Ϟ��+
�ittv��o��?�kHZ|_�K�^�j��u��Y$7��R�a�63	�2�fat�A�{�gm������r%jv�`��nRun�1Ӭ��q�7�F:��{�Ƿa˶Mx�ɧ�;�����݆d���;'hp��)��#a._K��� *S�$nz�f�J^+$�*�S�X��߼�4�#��k�����F1=�C�dbxh��}8��1�tL}�p��~�����)�S���3�lۯ��t� �n� �ܵ��q����uY�0�#Y���
��Gg���c�L�>,ʽ����
H�4�(�l` c�"ڻ��s/��&���`S�<��R|)X����?�H2bU&&G��׉L[�j�L�R��p��[�'s��'�j�t
�
4[r�De�BKpٳg���/�%Z�Κ��NW*Ш�\ǟK�>�2�17^)�l%������=�D��J5k������vdp������t1`ǎ~�����#�QI ���I�8,���� A%E��R�E��N<�p؍"��6�}�q�m�@��r^���V����۫�惬�d5z�ok��=��[sP�T#קͽ	˩C�	��ը;�# h�H��y�h� �_EW?���#�ƽ?B��l'��eم*HhT�^�l��$��չ��Fo�A�{���۱bq/k��%g�}	d����$4Gz��p�+n�}�r%带�0���uP�5*d������dM�E��R�j
9T9�~���,(�$�5�d����L
�����Q���cz����:|W�	h ;��-�q����pV�@uaZ5�	s[;Y��&4	�uC[7���>�3?�6�LmF,)�V������E�to�{�9<��?��Ǿ�l�.4�8��_p���G�k�P^��>w�������d��]��
�v�7>�q��ӓ[p�ч�����M��3��(K����'&X����������{�WĺM��ܕ�b��D�P�%���J�m���b�r�ž��/��zTu ���^͆��t�희U��*i�E�>Ar@Q�=�3��1����p�HY�#@�ϖl����ijf����Y�Lu�:z?�*�'�x^n��2dӀ�h`���X��t����{���k�X�]	@?�}�4~����G�En����.(zV ���1��T���=I���ʀ]ƽߺ1��#�?���[������BOO��Q����ϯ{	?��o��S/��t$S�}f��sC6hI��QcJ�z~�����:�h�gO���3���܌�y�P�Y���H%��R���Z.
�"��҈&�&�e��,�ڂ�?�!\r�ɜN<]���.�$!k�6ٜ)0a
Scl�δ������@����&�&^�!4 ��;� ����.,\��L�����fhN�STz"/H��5d:��;oT]�Qa�T�m�V\č�1��f��,�aNN��!�.@�LqS�܊��-d�:��o�����)�<N3��UE�HI�"vlF&��/�>�V���b`�B�B������l�1�`@S���W�ٶ_ջ������k�Y�θ�����g���^у+/>��8��k��1�T&�g��֯��I��5�X����#�։��
&�M|���1�kB����X��)�U��Y!�A���=!-=�����;��pswwW/-I�� ä�]+Q����P���E�.(bUR�9�ɵ�]MP�́����Hc3��=�gY� *�t"����c&?�w��@|zՇ�%$cF�G0<6�T���8���eՒ����Z����������1tw,C*��]G�+F�z�G&zL�1e�[B��Y�ƞ��q������U����$9�&�Jr�d�n��K��G��??����a�<%3���|hz�7jr��Y�a�u��A�d
��8�t�n��%��V��L;���?�b=	A!�35�7159Π�~�l.��$4C����ْO��z��6�i�p����AW��B�^p�5
ZL���0E: [vC�7�kpp9,J5Vڠ�ɀQ�ڈ�ĳ�Qf�D͖/B2b�U冋�K���� K&G7��m�.����Rƍ��k��[��2�m�RHj����pq���n�8�ƴ�N"�]#��oB��ù:�=�����0�}n���8��VG�^D�VD,���4����������5O����,.��.�: ��=�@~27�м"wҹ��������>^�8��޾q����l"cX�₏"�f0�Ӊ�l�#x������B>�q�|8��[���G iY���JjW�kg�%�}B Њ�g�Ph����ܩ���QU��4҉4�|�f�hooG�\GUi&B�1�A����Y�AZ
�D)����o�E��hQ#-Ϳ[��6��NX��
�kY��w�F��H ��$.:�$����Q/ѨՑI���(UG�l��;٣�&��O�����w�.W�(>��n8u	��@�Z�$��J�DUB?TlIe�~ U�s���I�>�PG`Y���D���M(Z����� O�Y���ڻ��RkBS��p"BJL��^"���zN�v��pV�ޏj=#ݎ{������A�-�c�+/�j���۲\�g�t��+M�d�Y��B�jW�k*܆�#޸/����U=�yq;>wՍp��瘔,xp���^��:�v�c�.+U�CP\��֣>�4t�ѷ8yچ�n+�W-`�ʃ!�IX����m(�>ϩ�ŧƑ�tcr�ƀF��s����D�g;���cgg'�� ��P�}����k�f��]�΢pJ���V\�ɏ�����*־�T]���$^X��5L�,�n+��tjX�b�� ���7x�?z�]�Ќ$34���Ys�W�n:w�{?�[��x%Vळ���-C�3t�Eal�9�]8t�e���/Ėm[�����o�} k2fr�x���d�nX���1�v�w���>�L�"�������gMI�nM�&�=Kp��ω  1-���XI����*�k��M�6�z
;�\�	\�tt�ó->�BM��J��T8�Me
��W3{}�/�pXq@�Ļ���䬡c�{籂H���Ai�$��;o��3"�F��,*U�/C�tZظq+~����uۑ��C6� q�����#&gP�֐I\P����F�6"`G�HȚ���W���J��N����!E���i2_�9�_�\Ʌ�ꆖl��(��Z���sxt�*��%S���[�Ʋ)�zӅp]**M��v�������ݠ���i�:!
�U�8l/-�(�z�j��I\U$�,�������U����̀����?�h�nx��*>*�m�� M�>=�W"���FC���QGyj����0I����B�؄���{�J�����!-�V�E�"��j�P��ȕ*X�l�,7~CC���zN$b�VˠJn�����Uy@�$]c.���x�l���D�A{&���!,��=�_	�<�@n@T\�j��G"���M97�:>p�)�)j��_���&t�-���O�05��/>s���J�L��oW`����8^��ȅw��g7��ݕE~jF��M_\-�������h����2otɶ,,G��\}��H���n�Hmf�"��H��� jZ�!ȡ|�0��n�,�U�=�M�c����!�bt���gS�2��c���~�K���Gadd}�)h*Yi��:j�r����h��X�p���'j���Uv������>���U��mˇm5�N�&'��}'��V}�j#c9��a;
%�-;��Lk֬	5)�
U1 Q�M�iD���eN�J� Nk-��1��9.�1fm=
��n52�}=��u,9p����dzp���?���wC�FK���+�TK���&''YPL,F@�Rn E2�YM��Iz�\w�y(�L ���u7܅���d{�P+p{����SS�q��SW�<� YЙM�%�u��8�����F�z��k:*u�U�iIP��99��13�Vi�ل��Bע�a��GI��
��aN��&T����	h�.t#� 14]��V�/�S#��ݯ0����EgG?�Ole��^{�����8�5tM�� ��s�7c���caSx=q!���Hr쐝�]X�3�499����G�7�۷#��@�d<��G��׍l&ӭ#���,UC�m ���Z���{))��1U~zW~�sI����t� s��5������w�^7�a��zV�b�8� t�QS��M�d3%�!��d��⺛v�v�p�8��T��p�vȾ�j�C��]Z��58x=�ڡ&��b�6��j5����v�\T�<���g����ϭ]��=����X�7��`*,��D�Ն@�e
�P�jLf���Q��*�$�J8�Q[���0TZM���p�����I�K?w-��c�gz�N�R��֞E,I���T
��.'�()����_�\���S���K<��[\�0=�'��P\x��\}�	|ዷ`��h�h�ة�ǲŃ�N%��_q��/Ϡ�w�V�j�u��<<���i���x��$Y� �FajV_�Q�넃a6�>��հ�v�;:Qup���d�' "öMč0��\�@����u�L�c����}
�7�y�u*�>}^�0�y��Q)��� �!�,��8�4$���� ]�.9������6����Mm�.6���	Иl�N�{1U0��2X�����<���0`A�W�@�k14=�]bnPC�2�㹶�~��!��c�'B�DlJ;��R3b�0s_Ӯvv"o�S� ]Q�]��'�^AV���s?]V�NH't8�:\�M���.*����Ř.;����P�0m��E,�aMW~zW���yU�s�ch殁Wd�s֗�e��.ir�i��G:���G�C\���)��P58���6����?<#م@��h���i���
�d"�Pt3����8/�u	�xI K �[FAuQ�S���6(OM�����d��ڲi�9Q���m��a�B�d:n�=q����,�����5��Cg@��W�d{&��rQ\�
=e��ן�׿r����>s镨[":��UL�J�'�a��:kj
;~�� ����PA {2@[���l�;\����v�x��8�������Ìec��}wݍ�>�q�rw,Y0�c!�I�;�������j[�r��Ԁf@`r`��#�P�D�
�L��ۯDo�̥���哸�K�B��Plڨ�EȚ��n p}`�gr-�Gh|����-g&�0Ds̑���3h�يn��k��kn�3�"��(�!�d�@ST[1��qN�}��E��7�N4�-蒇��u�r[`H\�z�|X.��%3�1<UE�} Kw_��/<��G��f�
_�B[�x4��%Ē*�
Ө5�X��~�
�@	K&	�J�p�F�Ȁ&
ud���Q.}��[�G!��B�M��<z�5���o���-��*3�m��}LKB�{��N��_�6*MR<O�j�q��Q|��O�U�"wӹ��14s����'�Ȟ�    IDAT~ï�N֏%-m8IE�M�Z�л*j�� I�3���:TDݎAK�ʵ�NO�5����"�:|O��#P��5Q����U��ƈš��HDKc�\.��I�7��,��:v��!�g�B{�o ���G�T��p2K��,���H��Y�u�4<q=@nr�;��8餣`������}�G�t�C�J�i��,!p����a����pTGI���H}eh$ux2���䷡�'��n�t�DΧ>ې1�`�6�a��%ڴw|�F�2"fJeW������q�?���an4�����#�E��h%�2�.�����Y���/މ�ߊ���(�.���r%E?U #S.�ѨU��+�&&�����ıG�*S�Vv]�ж)|��{���7!ۻ��	T�٢]����F�ǟALhB�Ej2��`t�&����5@q;�b@W�À��bhX*z�d&�-���T���yR�K�)�"5�ʍ
*�2��/\+�4����lΎ�!z�;g���ڱ���-�k�:����Ln�ް���:��4C�#7�Ě�6a�s�a*�,�=���cY�4���\�*u�a��W�F3w���
�14�����}�w�}�#/n/�=�l�C�
�%ԠY�@�R�"�U�H%�\�G_P�H�c:W�(��Y"���LUHdy�وݪ=����G� ۟['l�ޙ��jQn%�4���"�e���:;��	�u5Dx$��Z��yГ/�[q�T�12�Rv14F��0?$4��j�����q�I`� 
u��͛��$P����+���D�Tw���D�H�v<Ɗ�R9?��R��K8����&�����|.*�!|����G>t�:�?�W^{#��,�X
)-�j���1�&.��<�����y�6<��g���=���!���y\B�4�bK�H�1����*y,]؉��� ��}�[ I�(�t��,jn��BW=X���,�G�055��.Jԕ�L�xӛ���$1@)7�T�O�un���0]���ܰ�Ȥ1�d(��*�Z؎f�(n"�q�>9yJ߁�W�ؖg!׆�I<�ҹw!�:�u/���}1S)`l�ߡU(�3F�l������&W���"�1����3�!�Ѭ�*	��a�6t�����(Y:
d���觼�d,ˬ��+0�\������!6��tA�)Y�K�Q�בJ��p����aLSQ)�q�ŧ�N~㼰/a�5���
��Wa�_��<�ܛ��e��f
o�M^v��F,Ҡ�rc4(���'q*�&��Y1�X؄]k�X�K�5J@�����ś�l�JȐ�z��ү0s!��%������5��J�"�lHJ�f���n$��)�^k�C��e-�D��|�LPhx�@ȃ�	��KGQ�ED܅& ��-xۛ��W�z����6㳟����_����V��!(�V4~��O�����x��� X�D���4��k��,/膡����;��G���+��� ���+&?5���4���ۏ=
��[���v�`p)�Z�7�3��.!��92�E�czD������"�����\7��=0Sn�S,����s�/]St�Ϟ+1���,�m�`c��E��i'�	�}緸�+� ���
5=6Dh�$gϐn�p�_Gab왗 �UH�-1�GN�����dn}S���p&�
\�"�]ڂ�0�8��L�
��nC~��E�n��<�@�l�Y�k�t��h�6jr;�ǉs�T �!����#:��)J�&@e�uIt�#1|��cQ1�ȝ���@V$��U�u�cs�R�Z��I��e�d%�<qM��Z��3/�B=� !��;��[�Wa� ͫ���C����ߑs�J1.գ͛��wBV	\��k�mJ}U!�<�<���WP��À����b@v�o[�&�#�٣bQ^����G�W��4�b�shl�Qar/�1�G�w�}��[2B8z��0$�{B(�����C�ۈ q�a��P^�j���&p��/���-g)�W��3|��?E��El{6�sh4��ѱw���D$4�B�2�w�
&�R�'����N�Ϊzm��c��+�ckd�.]}-��K%%�UBg�ezH&S����Dn�])�oG�8��_�t�%��ۿ����ihFV�Z�ɽ��hI%���jq�\|�|ĞPe�>����X,Pt�=lGnϴ��c���G�Z��ʡ\+c��v�s%�nہ��yغm_���l�N&�=��(;G�bP���a±�hk�ah���[�xUHP�%ж�P�b�A��8pj������4��4��!)6e�,F�����]('0��ψ��PRxd;�L/���z��%�j�A���v���8<��52l�I[�-���n���|�F芢�_w�����Z*��A��m�.?;�@4�GcV�9 F�	U�O����zu�y����'�8h�5���
��Wg�_wG}��W��2��7�֍f�DLVỤ���>�iU�j'��FP���
��۸=��阬S���@�$��HĮ� !0�t�f�~I�2{1<-Io0���|P�
�S���X�]GMT�)��)�����P�0�0�i�
�HY�BS��-�l�32��Bg��x�&�1߼�:$t�\m��s�@�N���F�ZRs�8�|���b�v
�}�~h��"0C����N�a6s�}�^�p�Šƈ�{�}���X���qd���ئ��������dZL��ĥ�����'��������y�H-\�:1@� ��µ�hV&p�~�p�M�Q�)ÐcX��&<��Z̛7�Yd����2�"$"J5�$a��͸���bӦ�}��09U��DM�EWo/���c<lV���p��V��X�7f`VGP�XC���:d���ÑR;�ߘ���5нi�V��e�xu����7 ޶��߯c�_".5�t�d�r��G_��'и�@������������.���H{�ѵ�#�Hl��{�r�E������G6-m���Cτ��|]�k��*TU��q�$<�[�)��@(��,��Jiм����yx��睓��w��3�}t�p��x:ˡu�X�u3���B]Ԫ3��5��)��j �X;Sm4AO�P��bJ��t���=k��3�7%E�
y�%n�q]AH�s,{AڂБ2<�4NB`?��D@���m#�N�0�Ga�O�B�5�IE/b|$�FM",���H2IB��Þ+�΅.������{8���A��	�]��x\F��Mhh��R4#�"�qiä�S�
�3�-�"�R��G���U���+x��h������*d��P?�<"�I>6�	�e��ԙ8�M{���P|��s!��DH�ΰ��&+��� �
<s��(����Q+��e��|�b��.�<�L���*�����#����oBW�"x��B��|	�l��ӪC�S����#:���fI�����X���:WB[�
(��0C��di�@�����?"��Ŕ���kB7��z�����O���^�$$N#��M��*C2�Hgڡ'Ҩ7,4m`�=`q��nV )�|���7�u�2;�S]o�5Oc&�Σ.2j��U�N~�������DX-�Wk�<^��"��@}"��K�ǯ��q�p�i�;ޱ�
��^s+���yU���w�Ϻ�/�y�pj��v�F[2ѳ091]���)�(f*Wd�AԒPtr�Q�;Zap�t�`&�H��^fֈ)�:��[T|�� e6����ua�/�Z?�`��m, % ������d�0�%bpy�6[6�-��NDp��@Pv���R���4���/a�e��>�E�ےC����ވ���y��lBp�����'FL�1h��3G �)� 5E�m�{�[_�/m��3�G\@,����9�����x���-b�<�	�YE��q�٧���� ?���q�7~=�YV�X��C�9�E��:����t<�t�aX��rkB{{2
�	�X��\!�H`��!�t��4D1��Qm8hZ.3
*�
.�ǀ.%�"i>ovh����@c;g��N����P����8��$TP�X�fi;D� I$�u�7~۩rB�����o%��x���p�yǡ=���p�-_���{�b�$�0�+�o�ē=p��[�f�G�W��Ĭ&1Z��74L���s�0�O�-$1;]$�'�D!�FL���u��6�0%fa(�@��ġ)r�A�+\�I�`��PGV�PP��㙇���O^����O<w�G����7���\�����F�M9�ɨ'�7r8���pЁ�����f��"/�ߌ��G<�n��Ka:2���,��<
���w��kQ�-�f�~&Z]�ІN��_m�Q�R4��~n�X+I{�4��m"&d�MV �+_w憄5!Ә#�g`$�	e���j�e[C�0�Ez�ۓ�S�XQog��4M�1����qxL�-��(�.�^-��W�r�@I�!�~��������k��x�[���4֮Y��1�zÆ'xAgD�/f�H+������("�����՟9��&N;���]�̛En,��E*U$s�]C�>�L&�-��z��nK��$T*%lٴ#�c��s�)VQ�4��;�|�I��8��9��uI"J�<$E��-����F{��1 �{	As�hs%C�g9b=����D�����g�TGQ�ގU�~���5J&5�v緱t�!����	T��L<ə�kz<�x[/b�.�˗�,^�lo�v��!��w�w)H�L���� ���F�$�GQ_�nQm��R���ωES����e��m� �)P���Sx�ɗ�]Hv�"O"%U���,�	���􏯜�O�{oᯉO6w�&N�k�M���/�}�hȔ6�[kE(ng~�$,_܏��,���#f�F�-��7:p�=?�7��	����\��O�Q,����ٳw��Y�&bS"�Hx�9C���`�hj��nN"��s|���ؕA�oÞ)zb'�+kk�g��	C�Q�MJ�ey��!m�4���U
f(,��T�'U+�e�~m�.�$Y47�S����FiRv�߰r913D�	F��L�QaiyT#��|Ǉ��6��z��nj~�W� 2G��s�Sh�������G��$N�P=r� c[���K��`z�E�4c��P$���Q  �L6�*���<�#Kt�z��d�z��%F������l�(�*�4���T�@)��G�0S��E�P�MZ##��݇eW0>��5
C��4}4��PuHp��mLm
��6T��8��C9�޻�+x���Z|0|��]���<��GZ�a6�S�0��p��B���z"����&AQ�5֋�^X�A!�g�*c�hK�L��F-��7bܝ�=d��k���Ǯazz;d�s�aX��)-�A�`���1�gl�����?>	9�9�A��z�)f�TIF�^���14��;�k������{ͼ�N�ᙱBm?I���E�N�>�A��^(�ǡ�T�
�������0���m��P��7�����=t�_K���+�5�Q ��l�ȎL6�8s��"-�$r#�X���I<;��� �����}�S���Ho��#F'�҄��h�E�{ v�ʙ��������Jm�E?c[W����=�@�<��W�(2���'r1��p _�-!�A �:�^��94��{���P�T�Q���z��]��iP$%�r�0e�63+�
	�"�"�����!�r|�!�T-�O�������b�hMy#�iEtX�:������9��Ѵ�k1.U4b�@��
�������|��·�-�A$H�`	�Lr������=��X�"�0�.�{V��ƕȜ���`��?ì�#�������2*�"��� ���%p��v�>ʀ�Y(%Qo���h劅K�bg���a��Wq8��B�ª�P�E�X�=��.��{/����C
��$�i�(�3[��ߌ���xT
��H N�Yg0M�/-�F�����{������D�	$�]�:_t��x����'��;���� �;��ܧz�)��}x�x ��Mo��:g�zf�v`�~���y��'0pzzzP-���}�r�Ig� ξ�<�~F�̘2��ɜ����U"-K�!�h����`���_�,bR��D�N�/�,�2pf��B�u&H�@��V4͝�g�l�vE�cPe#�qm�.۶�=�$�z��oLNe|���r��h('� @n��ސ���=c14_�����V!p.N+�֌��,(,T�O��x'oG�T����p�3K$�v���T�o�$��B鷩TM�	��R�Ϣ�PEL
�D�o���0N�����dy�y#&��ĸ���}�隆 Js��RӮq���X-�+1G�r�h�%*�h4��@�H,2���C�fh�Z��
k̺���H�폪C@�CBm�0�4����b��x<� ��u4\H-E,;#����g���r�5$�r�s!IG�XB{� �vC�!@RS��~GpX��Buh!�P��kڴCP/�a�)]���H�����]%g����8�o��]��֮�����&�z�Ug��R�BO$�;�F2�ˮ�����P�]����R-��	��f����݂����`� ���$�'|�w�GFs�˲	�>�;n�
�����Չɉ<֯߄�Q�E�fR�����7C1HZ
�=�">�٫ѷ`oxR��GHoZ���l@1(���1(-Y�ß{y�eN"�'C�^KQ��	��W�1h�И�1�p�!5D���6C� �����EN�g��$kp=�)�HM����O��⺅+�x�ɋ�O��O���=�㠵����}5�+	���c4
3�͟�VHccӘ��M
�ֈN��%q)�J�0WG�t�*Ub��rh�A#j"�u4�V)(�CX�&:3��P�S؆N��[�n�����e����\b����Z��+�ڦ�P��wB�I���~�>o��Ui���\��,�j�蚿'�{��HPD1������N2��M.�t=��Fz��~r���럁�܆�j�i�ȴ�@P�Pnx��&�t��n_
˦Q�B�6>.2�Ek@�5�j<a!y8>m1lb��aֆ��l!3j��DZ���4��
��J8�I���+���0�֠�*r͈��C��kö�9�s��P�%9��'����e�I�{ͭ���s��UZ���a�����˕�-��p��+�����^Ƽy�P	�����/n�@o{��8���F�YF��A.^�*�Xu���W<�z;d-ϑAV�����G ��tc��4��hy�s[]K����:A!e����zЗy����CB��^��n��C�(��R����L&���sP(���:n$�):o��q��Z*8���FԺj��C��"��J6�P��"��=d1j=���qq&QҸ)4t����X�B�hDGz$���ֆr%�n�o�{��nBo�*���\X��"p �æ�V�y�\�	]��2�/������gB E�����(��q/�es_�4U�����Br���ǒl��(�h��O�O�������T{4�	\%=sɥ��Y�������lK@�½��#C�������P�ڂ��i�8K��3u$���=z������Y���y�Du[�(�� ���C�σ ���"�����#HZ)�3�(kC�3>�^aY�麤��4�oh�lT�Hڳi�[�,V��Q\p��(��L��Maf&�5ϭ�kuϽ�Aw�<�����]w}����-�ޱ���7d��0� �{ͭ���s��UZ���aO8��_�厭��������VL�mːL�����L�[7�X�s��������]���՗]���#۹������I~�'���~�=���ࡇ�t.ό=���OӦ�C"˨��n��;P(
����{�ڕ���p�P?ҫ��n��X�lx��bi�G�T"�XTB C��u���͆�Y��    IDAT�n[6�B�X�ƀ�sHF�G�e��g��1��Ӎc��ݲ����Ud	'-��R�?K�z��l�d@��lH��qkȴ˘��x��qMА
��@�:�fFB��{���BL�i�G�~#/��^/��&dzT5���	�q\�L-�!˰ :a�%3Id5'�5+ህ�/�*&�r��C�Bgq��:g�Geb�@0�PI��-d�r#/A�&�5�<���  ����hV*��>��Ϡ�#�c*E'6F�xQ�A<�'�z!e=���&���%Kt��f�@��a����j_��-@P�hؔ�0;#���+2[e	�݄������ �Ncx�R�
�R�f4T��EV�J�	|��Kq�q�ajl�B���ܴ�%G')�s��q,Z���id;���q|��������� �l���q���]�
i����
�J+0h^������n�����	fm�9�P|��S����bŲ�!o޼�}���Y\�x�<tdS(�Lc�}���dņ����W���ߠ�g9���x�,�Q��n��rX�l6n܈ɩi��Qf�W"@�b�P���]&��˒�i{l��������]K�j�VWR�B	� p,�+%h��l�����.R\��>���7��L�F5b��̦j`�P�L�hc5<ል�P��a�c��	�iȭzE�x�'�}���'j�)r$%�ksBy�F�ܬ7����d��>����p��oÂ��(NU7���@5�@a�uh	��ݸ����?��@�b��h�
0<p/r�����x>	�[#@�a�s�"M�?��G�'�N8�(�0���ܲ+�9�*kRKc$��"�!�ƃ�ň�H��,ph���2�э�#�:�зdm�`�tQ�!T1��O�)n�ȁ�Y��a;АJ/F,�;�X��6���&���E�2��	��LWG��ݑ�^�2e*d�����R� d��bR��̤خŚU�p��c`` ##c|.���Ǚe!&�1��m��I�M���[_	�^@�0��l���l;�s�^زi3�oߊ���&?�u�!������n�r�����MӞN:��y��y�����>���;!��o�g������q���d�Sp%\���۶wlwlvlg'۶m۶m��c�c��ϩ:O�u=�9��f����S�#��ipAT�����'�H"���m�a8n`�
�R��b���}��a@ȥ��*N=;���aY|���Y�ʲ�0��o�D���I�pK|���ml��N���C}�fW�]���o��i{8צ�4��U�����$M^���n�=����R�"K��<]7�O�
�w�N_�0!=Xu��amł0l��3�Pnrd�b#�������o�^�I)o-�6p��˄��󷰻&b���'�Rt���C��$�9@�ޛ��bÿ��n�HwBwHd�a������;�����������(���I�J��ɀ���Z�E���+��O8��6�˩�LL��7�߻�O:�ZD�E�/�+�Ԡr�B��T���@ 5�&��s�҅q�i��C1������Ӑ�i���AQ��{�7P���b��"�����и�	�h;_�J!Dq�6l�82$���a��1�h�)S(9d�
�n,](�$��` [�ys���*��d9g1{�_�Z,��8�Hu��(�s�����[�����K�5o�{�=l�;+��uqB�diڰ�������?��;؛�SiW$�I�K���=ߣO^�Y�K�O·������x���	+��R>u�I6�=����L����h������n���Ř�wt{��S�������������7y]�	"���=��,�,�a#�x-4xu���a4����v���UȦ1#�3�z�\�{A���ַ���YΌ�(kǖ�?2^V��Xe���w�7ӊ����k�F鸣Q����h4ov��pw�\�E6E���GQz����R�ׯ6�U+,U��<Z�%���0�aP[��M
p��N!��Yh&�b�x�Q�2�8J�?ubn4ܨq�����k�lԟT�G�~?�4;`�ysF�a
��cp�}H���#�W�Rѭb�|��H�c�1}o���R�l:��	�ix�i,t�a��1�\�
ft�9&:|n���
�!Ȳk��_��Q��V�(�k�+;`�ⓝ���m���[g9� �m�GrV��忉=���97�(݁���p�V��]��/V��;��.�@-���<wA9(��Z���m:��7-PJ�Amb�q�D	��T�E�C���_z]���)�j�����P��]hKp��ޏ��� O�FdsTr��6���#[�s���R�߀B"xmj�`�rTe�&�ϕH�� ��`�@��ȗ;}N^�}���>eX����2�:ZSm�p�3aW�{v�s������@ē���u�Q;��+�=7���D������{��ὲ�l��ӧl,�m�����(KI�k�ܼ��f&���S�����@�����ٙ�9��Bۨs��Atv� �f:./����j��r *]/�;F�'"��D.1Z��*:l$���'L�mc�"xր�UZ�:�k���&h������*`�t��ᆄ���|&&�c��&I@�Ch�+�o�K����&�)�^���[щ4Ԉ8> �l������f��xQ��Lʻ@��Ct�㷉+0{�r���g�v�+�KU>�@s+T[-t��2e
�����[���'i%a�t�g;�<�����?��&�1��r���$�QFM��#�S��7dl̋g>�m���l7��Vl�{=���7�o�[�W
שU���m�*_�ơ6ܟ�K8���U6Fh�h���
b���	��"uE�أR�#�U!	$�Έ�� Sn��*��Hy~'��6-�s��
8I��Uz"��S/J������.�FYȯ�O^ʎm�#��̾�CMU�s� u!� R�9�.[sj�?�}���b�\�=M_���]�&�4���L0���͊�Ȩ:	����r�U�t�|v+�5}����e��j)���<�����h%"pאk�ݶg�K�"�ͽ�M�4J곈}^h"l̷Nż�ѓgCG2!��E��_������rIC�^z-��4�H��_m��ۆ,Z��W��3CF;X���i�I����s@}}'0^АJC�](DlQM����]ۯ4Ga9��8<��k�Y�������a�i�-�R6$��9V�����\O�2�q$�a��/�_���'Ε�/�u2@B�S�b�	��`�#D:1�JNBsp��x�[!*3�$�I�p�hQ�	���x�q��Ǚ���X݂X��*[���Z�����e��`�_�i��̋q�2�z�vz~4Q�."1��d8^��I!�5 ��2�|=�����gM���Y��~���0�]Q�MOcL�o��9��5jm�0�a�+!�P�;Z�&ӄr�.�%�_q��م�cQ1��|֜�ҡ����ʈ�G��	*��0l�,�O�{&
�~�-Z��M%r[�g�cLgc��qy@��vp���� i������MG�Yh�e�c���E��#
���vU�a�Eg���E�@�͕���cМr	�G�u�գ��o��^L����#����WeeM��O��a~{Q���I�k����V�y߯���@�@�U` `X܋�3'O�&ͧ'�Ѥ���:I�nG9�u�Ʊ
�Qbv����ݵ}�X�_O�݆����� ل�W��>_l��
�r�%����[�\� x��X9XSa>�0��gI>>��.�ݒ�b��6 (�(t�V�{-.�DGHǏ	 Y��M��g$�c�ء�+

4D-mV�*�y'`�����=�x?~
����9zT\FF��W�oJ�D�,b��w!��"���X\Q�+�F��W7��/��EV��tҵ�IqdI�g�����w�ǐ��ޘ���bY,��V�J���5g��ڲ$�Ub+�=�8�v���x��w�4'i�lnƯ｢V���3��p�M�MrO�������)T��o'�n���q����v��r�@�O�-1.Rȶ]������u��7���;��$)�5��2i���ȴ��A̇q}r�$	����[���E�v�v�Q��>/��mHU�<"����W`�׌'[� �3��-^td]�)"��|�
zmA}g����R:���3�u���aE��bB�I
�_��X�&�x8��{7߯w��!?��G��<ɄCd�~��a�
�d$�P���Sd�� � ^��S���Y�8^$nx�O��tt���X���Eel!���#�{��a�	(w X;|�<v�,�(?�6��Q�i�Va��܎������A$�;��k��w7Iʼ�H�a�Kfu�Fx����7��5�H����?�~�-S����E�t���@9�M�|�:]��%�6���ƈ��#/����-<f߿�Uٳr�J���r.��ɡU�M,O�S4��C�>>��Ms�]�T��>|����g�r+b��^W�F4�A���[XX(�VWA�u�d5`p�U����(DkF:���F0��>�\$c�ks��,Ahw�x��8>:��A=�d�$+�]�	t�7�c�{^(0$���Ay���'�c %�AXb�g���}��^��Lr�PB�=_�E;ԍX|Nx�ާ�TZ�:��h��=b9�ݪ Ux���[lͅ��Z;���V�Ч";�&u 6�
'�0��Z9��;�Gط�[��tn 	��V��W*���/�����K�97��)	��'��v�x,�}ؖ�m]��o�@~�u�@^��(hj�-h�����<��<W8��#AJg�P���������$!�Ǽ2X�N��#����K��bʚ��*6ʴp`d`��D�?�������n�?�tHpH�vH���[�������$�c����L�
�Pg#ei���=��T#	����A��Ϻ�]���-���\.��@��;jN�u� /���1�F�WƆ�؀8�N��ٴ2��,Z<)x>'�r�F���#���Cz�V����M��1E�)�i=������%�H���Qwd����^��;�F߮��!9|��l;){�tV�MUa6�q�>��Б� eIC{��PJ�ˣ�q�!a���e�����2E0�&�Bz�8�$���]�Q����]	?_�;c��Q�h�>t*O�*����9u�$����ȥ��s�.`F[�Hq�8~���UJ-Va<�y獓�B ��x���ϊ���9-lmG{<�*a�"�*V�
cn�#iA��P�mTH;�0��c( �&���}��e��y�|��op�L��f���)�;�Z��4q�q6\qu�[�	!;,`�ӡ89j�H�v�˓�?�7�#�Wp�7[��wᐌ�C���b���1s���_y�^q��-e8x��/�U��)�������^�U*���b!/��ދ^���Vm%�3�u�a�Uݸ���chղH�d�`Ma3�6���O�d�91[���,��Z߳�%*|TLi��U�ӅQ�ps�yf��}9�V!�\�\#"Bd�nc��̋��}���[�\�����&�������C�_�g�dF�+Ы�p�׃�5Æ���e}mc�<�����)h����V.�0�Fx�-jot��`�^����ޞ��&���2��X�2�)ft8~�r�҉�jQ��u��fw14;@�K����&ڄ��P9�(��K:]W\�E�e۴Q�#���C��i";sV�<baЈܻP,I����9�9b5��@��հ���΢��[}�Iއ;�������"� �"˽������� ��qo��6��߽��O��\��\(��@�)��	�N�z9��I���W*I��2�U���!�"1{6��1��4�D����+�����ʌZ�倌�1xiq,|cD�v�^�L ߦx�,�@!Įu´K��ۅ}�k�q']u��;_���j3��@�M�!�/��I[F��7O�%�o$��E6�pR)R1���V�q3W�G$bl��kYW.l��Gh@�<�=�HV�d��|���,�>��ɉ'J��9()M�)0���e�VtL�lu�9+��ߪ��������Ik8�\�S%��O��`L�zrJ͝��ɄN�M���P#t�($��Fˠ��v*�ļ��	�7�K�a�%ʡ##o
em ����ܖ�
�s�ނ��&�����6	-K.��a+櫑��6�L�|=Â�u-~�P�A0�B7�$r�ﭽM���膵��Y�z���ZL,a�kkGT���n%�V�Q����ˈޕǏ�"�¶e����f����S��ҿ�8�ኘL/��� �mm���r�uı鿦\A�[E�r�E9̷��؊�{��x`w<�c�<����\����$��o�,M/��@,J����=�v��tt`��Ԍ�ø�~�>y,�$'��p�r�M��e�W0�q�!�]�=�ɜ����K5��yj)˴c[���	��q[����ӕE�Z3��L���h�X�� ��0��a�vR䀧�,rx��gg;��Q��c��R�J"R?v�`���)�)��>B�wM���i�Nۍ]"X�I.t�C�PY��MV�_
�?Ƶ=�;ؐ��:���7�P���9�5���!��~�_�n{G>�_|������w�G�7G(���v��k�s)j � M����S�
'h6
�D�ϴ�Rւ%�?Y��B��-Vр8���H�����N�GX�+�r�墹LN�&�\����ζ�H�Wm�YV�7LK
��>n��qa��Sw�9R������6���r{ln�$�d>�bi�F'�3�-1���얮�bq6�&��`��e�K��6-���7!���ت�!*��Q�`ͨӝ�:G�;��LYR��T`��ܻM`$~г���Gm�L�#����p��'(�&���",��e`�=Ml��3��=�Mh�j�A�lT!���&�^���l�J��V�0�`TL}! "BQ]L	"�	����`�c�d2��3�-L�U�ZIߋw^�u�KHiL<qy~u�V�4%RT	�������Ty�	Gi�0�q�dI�&�ĉ���1���$��B��.B�K�WCc�Ĥ߮��z@In�X�=V��`��/7o8��V�>B���2��q���6dH�"����S���j���h!q=�zq��Ks�W�|��קq���;�S��]��6t5�oist�b5d��W)�ȏ����'jƃ�z+�	�љ��=H����(���Ⱦ5� �:�ﶳaa]��������w��V�`?Kjғh;��4V{˟}�kuK�\��.D(�?r�nLC��>Ռ��j�����{Ma��I�nV P�D�0�3���B@�<.(���]��$C���]�GSgNl}���Q�X���g�?��$�$u�������k@�t��\0�� ƪ])<�B���e���U���y����87��BP�D6��O6c 6�FL�w^�����D�����"5�Dm�<�>�lG�l��}�r�b�	"�Z������z󜖩gE�(�+n�{�B2�.�߮���@�?��rne���u�%&�^�f���&v4��LR�B��q�0K�!�Lg�H��f
���4Y�`⾭N:���c4{��P�KȆ��K�C�p��u�V@�n��]�c�k�f���)0$����t�L|XԐ����5p��2�q�U����~�m.*�;>ͩ�U-�sR:���M��������=�n!Y�b�� ��ڈ��~����`���F�R[�ܭ+>�6뀌�f'>��,"~e�
�� ����B��Ua������i	�#At����g"��^h�����^b]�0���c��Ң=�����0�r��MS���2����$v�հ}#��%��C���NEX�äT�����z*�$u<^a8��}��N����w��1��IS9I��j�xL�`Y�GN��}"���х�]!�1/#S ��1����	�K��#;���$bLt��A�A瑶̮�S�s�����\Y̷ycw4Vz�<�/׆ɝ7a��RJ@8���"�4��@y!fTTw��@:�/r�[7�ȘNq����"ݦW�+q�]���^��.�2,�3�hP(��$�q@�c�%�f����D]giȲ�[볲��*O�L�vqWKT˛�ʣ:�`��Ť5��$���x@}x�SZ]��(��WƳ�$��������'���,6�=k�����L�a���+7��M�����!"��Rk��tZ[u��T��o�h�L}s�m�␆����o��kt�V�O!è��n��xa�/ě[a�af�!%��X>�ֻ-�~Y�Vѻo���@�'|���L���y��F��Bj#�\$���-�7�M����X��=7�E+�hS�N̠��_F�c���D��]9��-%#���"�º1���t5�3�c��y�^�T��N�;]ۦ�Z�7��bD�g{�x��i���
���N��zVW�����a��Q���!_�0J"��aT�}XX��]1}��-R8�W@���"$^��j+�a#~����s�P�����ҰÁ�J��A��_<Cp�G=�S[�����I*���})9a�B'�U'P��/
�r ����/�>[Q�l��C��R-y9��ּ)V�0J��A�hH�s�V_Rb���&=U�wI���yj4,����z~����TJK$=}X�:6����P	��0��Ii��U5�������-��;�A��1�G5ȇ�U����a}��6h� �]5sv��j=�σǄ�ܙ��A���^��'�����K�������`�΃�gqG�e��Qq��h�6���yd
���kРqs������]��7���S�ª��®��݃���B���F8���z2�ӊ�e#��o)��8��t������_]���\��E����މ _�v)C�C�=�s��@�y���=2:�1?m �����*n��ڋ�qb�m��(��8�X�d	ku�l./��f9i�({�%�,���o����~�;����S������1��5��G����u��I?6.Qp@=t� �2Q�@QG�~����������%¬*W Δ-$�2���k�@����� �S��%{������l(��c5�@'}Y��`i�DD0i�r��N�>
d|��wG���������I�*�E���6�g.v��ۙ������g������\Ҋ�|T<񜔧�2������jHЈ �F�R�?���/6���cvU���R�������S�x�L^�4ET�v\��6�׿	�\���,�>����z��&|:���N�B٭K)�|<6#<%�dA��m�0��d���d���]n^��Ͼ�ː����D�Bk���M��7�#q��G�Z{�x�M���|f�d[ܨ�hu}'D&� ʚJÏT��V��G����`��n]8���+?\��u@����y~���?d)ٔ���~�5JҟN�A��r�Σ+O�f\���!�eV� ��3�n��&��������BѢ�'�eVw��o��Ah� :4\Տj�LT���؜�}j��p��TK�,�on�!���T3��"[����Re�6t\t3�hJ�D���X��eB��$F�&�CbcV�=F��T�v	�8�i�C7?�`x@�q�Dj��L��__\�`���ta]y�tyy,,gn4�~27�x���Ȫu1����9u�CHg�"�����ȍ[]��b�<2:BL�ψw�%P>8�"��h;.*g`J�Xw�D���y�XF�J�y��~)4ὙJ�2��#����t� �!�6����'�� �r��x�$z�Jy]���t:��1~��4,4�'�U��O��a^�q�~[X�qo��b{]!�����Q�g�~v���0Y`��C����p�� c�?b8�?��4;���C�u=����؄[�x�q۪�Z7tEӛ �cۀ���5y�bgϛ���G�ٶ�k��f��B��� 鈯5��(�+f��&�b���5SpT��A 'qB�<DzҠ���%�@�����E��u��P���!�E�.��-�Q�5�BÎ:�4F�$N4�뵆���qdb-�=���.���~@�h�{z�β�a�Ϗ��YJ�+�n�r攈�I/3�D��<��~�A�8 cd���Y��T�I:�Km�,�å��J�����x����&�������㰳&r��&5���`+��A�,RA�\qݺ�T���t����H�v��'`��u�x�9>�j��rbǋz��i0�����9}�4��œ��.�!��?N5v.&u�Z��g��A4�!�<]�N�m�˥��/�h��]hڛ����A��RAx5)�2����+��n�Т��^'H�k��ڰ.��΅���2\.&(R'ʁP��'����IU�#~�C��{"l�R�B��,���̺w/��}un��?8��m��T���rT��Y�5�O��^;L��1�(Q��y�Y��yzb�B�@'ep8��1��ssFUۏ~w��T@I����Y��k"�g��"Lr����k	�.�c�ܭ V������؞�?����)�d��h�ƨ7Y0�4@��+P-��D:�;���kh���^�S��S!&����Fr���K�Ѳ�"���I���������e[8��X��cT?� �� ���0����_�o�~�d6X�����m��R��ߵ9�ma2�K�}��v{� �k�L��J4RQ�Դ8� � ��4}1B�$�}gK��h^����=��k���_�W�q���ߌ}�^��Y��Y���
��wY�?�I�n0p����4�=����vww��Ҍ��$���jr��[�Z�
v�V�fN_���`k�XY
�{���pP}0��d�%��6MiE��=����R���~��Ƒ���rl7�����,,���<?��oWj�ZVF�H��΁�uI��X&^���`d�>�����1B3t\���O�����(qz���������Ѣ����U���Zꄝ`�V�-7I���a�ڭ�x�A��ݽ��0j�׃��R��Uj����"S����Ҏ��lT뜈�Bn�����H�MD�~��ϻ� �r�|�Տ
'L�%�75S�����?As�H"�`�Qf��HO.��.=�T��F������9L�M���Z�:�C�J�Ƞ8LQ����YQ����q�W�2�3tV;��>�@�¾�*/oJ��"�tΦ�!��`�
# U}����cC�G��a���t���S�Tfl�,���8�iV�h鮡ʋr퐅��ݠle�a����@��_���Đb�Y'7�0)�G1����V�A7��:�+ g,hu��0�v.����b��'�yצ%���s)YM���<��m����@��rhBڹ�uRHe�TN�yq�#��5X�<b���l%HǏ��-t�l�'��V劊�1�a��x5��B�!zܠ�/Wu��jH�W�,�A;��:��b�U�v�?N��pE���i~��±�ג�]Og�2FյeFӵ4��"�D��u�E�݋<&�;�`My������M�u�[������_E��@�	��v�FU�����m��O^dsG�B|!YI8���¾><�\�)h|S 64j44�ɣ�#��z���hz��rH=��ٜD@��n �>΢_>vb5,��SDC�<Le�4U��c�tt�h݆���E;��s¨n�00ֱ{�qH�
�m�֬Etm�*�Ml������Q�P�W��Ȗ�[��PW")�>�[Q1Z��G��2��^ߛ� /7��Yçd	l�hql�4gH�*HБd�u��I�ZTQfŅt4#!�ܬc�U1R���t�:�8�Ɩ5�%d�	h�w��.�r˔!%%2!�S'���{�2n���\ɘ%}]��}��F��J�ѳ�~��l|i���bʁ.�'��}} *f{�����ӣ��&!=y��Q�fq�'ҽ�}���R��C?��h4�?���z|w
�65�+����̞BV��
�	P5�0@�����{/,ݱ��U��E�n��r��5��~�<��	����b�X,^�O�z��t@SR�!D5�uB{B�����8��?���'�c�ç�����,���l4;LJQh�N�O��v*�z�ݹLg�y2{��{��W�ic��܋�m��E��!y��r�`�ձ�i�8��z�
�
b�ˏ���iı���"��~��<�+�|.�N=���+�]�b�`�"�R_�3'��b��+���BX�2�=q�);X���}<W�.�%�N�����f�����]1�T ���-�_�F���{)�dO
�&|H�0Z�����"B+��8�؀��8���3cD9Sۗ�^U�?��&6�����1Z�����?��[J���H3�H�cB��P�Xb�;W6d�~��0[pDE��Lt����7"��!�^^_K��sD��������s��;�}��I ��'�$�$'l�_\Ȉ㣡O����8��94�:}����D�r�U}x�<?�5�0��z7�mx0�c����r�($���1�W�+�+xG
D�v�DB�/h�5*�*��A���h��I�Zތ#��&UG�Ѭ^��b�����/�f�]�}=GNV�x.�ib����*�4	8J��;4E�!����c0�"l�m;Sv�Wv��H�;>?���}0~��77�R���o������n�[�ة��w���~?h⥸�PWc�d�t%E���j���P�m�j*�V��V\K�>׍_g����U��9��a��`�|�j|i��R�)����5���ڰ0����NhF[ �2�7����t5-z<W�Uh����u8����V�W�H{�ؑ�_B�m6+C~P���G��M{_��ދ�#E�V�g����M�z�U�*��5��_�<��5*c"�)K�A�N
[ס���q�v)!����ܘ�Z���"r���)P�UGk��t�t�jB ,�N�=W���6��Bx�Ǥ*mI�cL�O�OG�ΐ)��ʺ��E�[Cf)#�/t���������a�-AM�����3�	���s)H7����Ă���'R?�q..�eQ�v6f!C��O?S;����,b���u-;<H2����K)���ق �@�Q+2�Aнj�'#�G��׺��v#&
@LO��}#��1+T��0�z8os�Ѿ@{��"��E2����^1�z���;O5x�>���R�jC[1Q>�;<�l/N�4$�U�_����du��Z�����lT�����p��7q��CO�p�����<�FӍR�`_{��Q,_!ʉb�Z�s��jt�6�����Ù��G�F��,&��#��f��YP[t�S2yH��[���`������������7�e6"~X��_��s�@�0"�bj>��q
��Xm⧽�&�O_��v�JS��H�wµ�!VZ9���[�t�d!q嚝�)X�&:��P�F�Qh�a��,]a��ʇ\\�s5T�)�m�D�k�zBA��� h��n `���U\�Ҏ���I�߼Y�g��]�T��{!W,L2U	�Lz\�MG�4�b�<�DudRl_�7�'	�BEě�G��x�8���Io&�q<�����a��&�~��(�שD��xZ��]pD��y����q^��h����?�潸�R�)Z*���{ݲܰ�-S��oF�n4Zp�ju�as�q�+�qqi�2 F��*e�2? ��ik�ÌP��n��9#����[���7P��;�&n=�H?��1C�����X� 
�iFR�D����Jf��r�n0?�
	r�Æ�� %O��@�;���������l�{΁�G�����_����!qָ6�8֪�Ww�>�m6�GC*����Ed���p��:�"�1�b@�)�� lF
j�:0|���5O���vl2��( ќ`?��1_OxȐ[2�f���/��8�%b.�T�6c8�J[�P+(�z�/���_�{R�<�kځ	����;�7�&V��@�8��iၡ~�| ���ů�Ur�?����{�$2�B(�XM(�5��nd�T�/�ֆ�d���������g������I�!�,H����6���	��?�ӝu�~�K�,���L���p�7���>q~���U7��?񋐩I�&��?�Lp��������}Tgx�o2�0�RP���]�^q��J��|�L���/�����2�YE;`ů��Љh�B6���@��������y^P�ٙ�L�NXYs|����q/I{���X��YX���f:�x�F̇X	��F�#����(V���-`.�F��K��O�JrjA���E�^'
��7�3?�[ R�d�fa�w�D���aJb��='�������i�zc!Q�e���Yw��ߗ���Q6��Q6��o=�M躪)�m����k[�RY��\��y����c �&�.���f>���}o���T�"8���;�c!�~�a��԰&Jx��7/�`/V��su,7P�����`v���|D��Qf���k�Mn����/����<8�+�vN0���q�!�e�P*Ja����'fu��b�9z���#\n��>����Jň9k�-)� ��d���.�!�=ɐ&
��䱅�U��x#� s�<�r�%�1�Je	O�Z��,bzJ�,�#g��8�Ϭ���}�Q����H�QήI�,�����k)'����'����g�". �?���h�E%���П�WE�1��RR�
1$�H2�4�w^�-�j�i>�'��:���'����%�H��*c�QʽMX˙�K��&񨦆�_Κ]GGG<D�=�5O(��U� �����0��������ެ�m����'r'�$+SΦڟB��7�>]O���{ڰ}���c�j@�v��L(��/S
=���:��������16q�s�BԴ�L��jM��`/;|>g���;f }�]X+�ElO�W
�?.6���{�W����ց��w:���/���㬟��{�x��{���m��O�v�hX�F	�/5�}���o"�ÍK�*�է���P]�0���L��nX�DQ<�C��N�FWBIXD�9Vi�K�IpKZ��qy�#���d�ѩ��F(�(� UG�A��|O#^'� Nh�w�TC�^�]��dtxb�T�����OLmJ�6l�F�a�F�ٚF�@(+��)��"Rupzo�I]�s�$(��i?�+�cf-`���訉��5�w�"v��vA��g>3�j^�Wb ���ʞ�+}�� #�
Nɻ�َ���Ͽ�����ٺ���Фd����a՟�L[O� %��I��|n�j��L�IMp�}9��k��K��>��Mψȣ��9>���^1�?�z��4+�0X,�A 8y0�jy��!NHRp��d�ڱ��A�G�� b[,Ӡ�����������3����;g�-f�s�};;�M�� �pz�`�8=�3�s蠎��;(���}M�Hf�Ll��]�]Xn�7�d��N��S�
j���8��=vms���=>b�6�����u��J��r��l1be�s���N��ZS�����?玻�3�4�����󐕚Ye�3W���>}fmw�F+��q� �eVTX��g௕�����HΞ�(�g� ?�\ٻ��	���;��L�#Dq�b
����1�}����<�xd6����6�
a���lR��a*<�Ru+�����uiޡ������B�{ŭ�qr#ϕ�'k�Ȏ��wD�|�*�Ԣ
�;��-D@�*��r率�$,c�$s�iL� V�m):�e�3M]U�{���s�C�'5�U���a�O�h���7��&Η�E���Ѓ�i�w�S�0Ɯ��h?&O�0ܬ<��1���!L�����m���\%rסގ��8d�z�o�m[aT��.����G�Ƅ�Ϋ��[�j���F|�<��c���2*�e~9lN���m`�S�f�#�6�$A�ë��i���/+�ğ���~�N�'N��^�OP����8���u�8�}��S���$m\&������F�RK�.Sy��Rb����;�L����m�o�[˃̈���	���u�O��B�M���1���I���o}����<) ˱CU��Q�0���(�:�r�G����t�c}�	܎*,�Si䂌� Σ�XI9k� �p�靆B�4&)��eS�t�_��!2���"�j�XQ��Xx̹~���������&�[H��v셏�����G����;o߻f�S"Gt�?����Gg�L%�i�R�I���)�����Kذ�	Jvt��u'�t	����8v1hQ�f�'���am3�|�1,HB�WJ���Xg��g��@����_@��l�Y[77��"��i�I<ᒂ�ęlg"8^K'F�Lg6>ι��ķC6a���3B���:i�3:����oT`��sT�~��F��}�� ���&Z"���+q��@�j��T�Z-] ����¤5y�t\;�1)�pʫ��ٿ�+g3�܄��c���t�&Y�ċ�����V�Jf�K!�Ŷ�|lJ=nEN��)z�N�}F���zܮ��Z��akؚ@�0"�}	b��k5��Rb@t�9��˪�ixaydJۭo��͍�{�����4R�j4���E��-�g�����an@��/�O�д2��Q�����U�����|��..<�Q��Ĺ�KdqkRދ���jj|^�ۙ���	������ˬpWd��sg���i\���Ie�7gB,�ĥ�x��~�� ��ӻ���Z(�e3���RV��ߟZ=GU\D��P�ގ0H*E�(����pa:nvj�Z���l��պa�]�b�G�����ZŢ��zAo�`dԤ}�Y�]�ykۋ�wo]�����TD�Q�&�Wr���R� ���GYD�S�+VX1&��o}�$]�D����
����
G��m#m�Y�M�M3T㐸�%7�{{���Xn�ﹲ6���h��j*U�܍��G���	��c��TT�����L������X�3E��:*����2d�R�п��8���1*|mQ��{m�#kt����NN]��t�����d���U�(⿛��4;�Q���f�������k��i�>]؛O屲���͜��C��B����x��V°�)n#��D]w����N�,�vVT+��zb� gV���HصM�48Qy���lo ����馾He��V9Ǭǜ�'�������(x��{,t�Ev�M�ĕ��1��z����Pǭ�z� e@���a��wt�1�XWO���������VVi��y=@����Qu!�S�*~
t:���];_"���R��̀?���B/d�=7\N�)~6���y�������Xv=��/����Á�^B����K�C�H�5�4�m��y$�Hx�:(��BJk�r�`%K E�>�8�&l6-M�x��b��Sp�m��&̙�^{����〃�ᨣ�E0�������+���P�'㦉�&��CŖSƁx�˥I<��CX��M�j&��<x�\�������¼��cԨr`��+PSۀ���7���ے�Q[׈\VGA7$0�.����t�[l1	4�캥�u�y���o�08�w�>/��
���_��:_,��:�$��θ��1u��p��!�	��חŗ_-ë~+W�ǈc���#;���}��������F��7\5~3�q�͹n�8������K��ͷ��gK%qx��v�y��*��59
~��W���pɌK��}��/ ���f]1+׬����FcS���?&�_�z�֭CsK#.�qjk�2Rjo���_/�g�-ƻ����Fv�����o��0�5�G	����2j��#b�'CE0'�+,�`D�'��1,�F1@�_�zH����W	�s���Bpd2iR�A�B�=i�RG��_>� U���s�0_H Ǉ���@k�gJ&��z_0(�8�+�3�����EҤ8�*�WSS�حW�Y��c&��O��!_H�0��� -�]�%�We�����/,bo�#�"�ҋ&ݍƦ�FN��`�Sx큋�㏠�]���a@�#��߇C<�[�Y�(M�bHz�Zȫ:[�+z�DR㧠ߋ��^�ҵC�2sJ /�Ml¦3��o���?s֙'���c�:��H���Ӆ���b�o�#Z�q�U�"�Kcǝw����{~���n��أpÜ3p���/�'F���f�Z�O8��0�}bo5�	>t%��%|��xt�\���
<���0��G���
7\�8���Fj��ꨯ��V2��b�?�s7\|�/��?~�O?]�Q�[p��@o_7f^:�'O������|��� Vۀt6��W_���C<͸ �L���+>�h�~~}�9���8㌙H�
�d<�c�F�x���x�ͥ�����4,\�P�O~���p��Y�{�m�쳯��w�Ǵ��ᰟ�n�=�|�)<�`6�8
���ht��Eo���K�mz�����������(���g������.<
{m	���;�B����A�1����r
�:c���X��-z��;&�qιs�b�*L�:���%��'_a����;n/|��:\3�:�Դ���U�-���ő�
��#Y7��
�c"���k�<�n�RL�T�WL6��M���2`o���CV��a;Lp��X��U8�EJa)�͊�1�h}=����T9��'�#V˻�7^�"�n��h�/ElM]�<d����N`L`d�Tz5�������¨��9����&pa>��p�bZ�,��+5gP ��d	l�Z����{b���fx~�g`��x�����w���932��c�ŭ�����r�H��vT�b�!��"�zō�3(�S���,���Q�E!����m.��{�68��3�r�h�04-&��~ ���$�{�}x���Q���>{탞�6����̻ÉsϞ	Ө�S�aܤhh���˖�%�j�K�bۭ6ü{.Ƶ7<���W`�sq�������p�z9��]���6\r�L���5���0<���"�� T�`�3O=���J���������ӆi��w��k�}���_�w��,^z��ꚰ�cn�~&��a�=�0\x�9���N8��3Q55t���y����+N����7���u<�zn͉��6�玘}�x��Ǒ.�p��⚫o���0��˰���C�COoZ�5�W_�_x��<O>z?��N>�\D���D�n}C+�Q������[oᢋ�C,Z�ǩ�\n?N<�x�t�>8�s�f]�hO�o̿�r\<c&O����3~�˓a8cH$p�A�a�=W��;���?�W^|A�_�v�N3`�=v�C.��[���/����1�v��� b��pC�W��U_��׮�� A�L���/�]gՃ%������(ѵ�IРM�V�S����,L��QB��5��	�D�U���f��eJGj�y�j�R�!7�K@�;9���D�CP�^U�d:+��^"Xf��X����c���E��n^,�Qț�L�+���9�e+�pq��K�rW7��ۿ�,�?�P�����30h�o���������c"�VW*B��d]�m���R6�B:������|K���(���$O�*c��(��p�%����NB�}-f\p���.��ko��[���;���'�M�\����;�`-��ś�O�Z�c�m������9����u;�&R(�!T�O�y���w�ô}w�uם��W�C��Ux��{0�;��ף�y4V�^��;���/���XL�i/�x�9��H$Q[�C:�S��kg_�+����:P[یR�u
]�ϭX����a<�ܭ�{�x��w1b�8��.�̙�`�m���S���?S��g�q�h]Z�8�C1v�x�y���p��+p8��>���p�;��.@8��H�W$�炳��^{���J�*Foނ�v��ξ=����DC���@0��d�N/��7�z�?|�d�<��e�?	�rQ���z�Cr�4\0�\r�l|�M���8�P�s�!8��w`���q�!?ŉ���@�XBA8m{�z�a��;��ֆG���0o���n6EƐ�Ry�d�r֯�ƨQ�P�PD
F5V�Bѯ�"W%�OˁFm�����OV��4^+ח��Q0����ٮ)pT�����긲���<z=>��o@M4 �VA����^'èJxL"5$A�~F��M2}�7�m�(ѳ3UhZ �|^�����YB,Vu���K��cp�E�I�ǃҋ�I�Q�A4IY=�ۀí*D*��1��`ͅr��'�4��O������0��7�'g`�c�\�ʹ��Is���,�~'�B�d?<(c̈&\q�ttw�a�3���o������ஔ�$1�(���)'�3�8Tڋ��b5-��ob���}�݌���쳮BGg�p͋�/�kW`ｷ��W]�;n�ｿ�@|�R�.�E��:�.=ntw��6SFa�C�p�����u,�77�t/^����M�f�q�Y'����ĥ�݊���	j�F#�o�I�5rH�6��}��us��Ϗ�֯�����ӳUG/Y�[��x�ᅘ=�J<�����>���\�s��{�=;�g8����a��?��1��v�V,Y�Wͺ0���q�v�����v�ccP���R���w^���<�O��*�̜q:��o*6�7�Le�4�����.��%��{��n�MEg�KUL�����S���90�<�n�˵wf�S�{��[�pތKp?ǅ����N��~1��9<����˟���g���N�����ƚ��}&b��N<x߽x�����f��K.�}�5�f���W�9���N���njQ�R���RZnug1`Qz����!'����CY����د���͠Vg�RAxRK��H��uٟt&�HHC(��/�?/��<;����w�l�z��
��8��z����1Y �E��o�5L��!�$xbIe��:5c�Z�{{�&��
:�Mp"#[&P��M(������Y{�r _b�H\�B4�9`�5����E���c�|gg`�|g��ǵៜ|��t�9�L�ᮖ�"�삻�ô}���M�i���ϥ�����_�����],[݉#'��	![,K���A�4�����q�ѻ���Ē�PS3��)�4��?��l�z�p8}���H�'���(Ξpȉ�~;�<�����)��sa��������q��u8�Jtb��c1��Kp���Ѷ��=wܶ ���C�;����o���9�,[Ӊ��	H%��NFy ;n7��z!�\��x�}�=m�����#?�����>�>|#��O��c/�e�$�p�]7�1R�c�:��r��z.�q��:p�M� ��W�^�Bޅw���:M��Ͻ��w?
��-��:v�i[�C!��ևX�УЋ9�8����8�̙����W�ig�
�N���|"f�6��r�s�U��o�
j6�J>���p��]w�<x�A4�¢��f�
��ȃq���������h���^���*X+ԧ�r��� '�z
F���s�EWOM;�n=�_�[���稫!��3��7�i\z�M�+$����&T,��`갪�jD'�P�CiOTS�ʩ!رu/C�c�KL�'���7���(�1�@���\C*��R����=uԡx�?b�}��G.ƺu�0+�����et�ͽ"����+�� �!U�M],�Q�!���e�
�{���Q@��Ƥ�7�m���d�3o�үѓH�/�A˘͐*T�+:`:��׉~��0�0�ܻ�_�q}������������ç�5�zp��^����ㄣ��c[$P-_�J�����@��,x���UԵ�AM�(t�q\E��͇r��D�:̹z:�;`K�{�EHDP����<�)x\y<��<��һ�{�FcGcx����]8�����c�a��Z�s�Ltv%P��������+�ą�=����6;]��N�ᖛ/������5+�Н�q��=����Dcc�=s?�;�p�y��"�1	4�6V�|!�\���̽�Z _9�j$LL.����5������K/����)�]߅_�y2�Z�D������kq�����1~�\sս��������3��'q��W��q";�(��>��|������p�!?�/q[��ᇯ­���;o���w>p/��3�n�z��E\w�s��8�Sq��	7���FM��l
��Nhin�#މ�����S�F,� �Kt��Jy�;�L��q�շ���@S���&�/�Z�s�>�N��/� ���"���G���ɧ���xO<v��L�~5`zE;fl+�y����_�ȂQS7Rr[h�SJXZ�n�JR90�(�G�	GP6338:��eD��ft<�����娥Qc-0X��Q�� �1Xf�����lh[�ښ �BA�#�p(���aL��d�E�&��E����SN.�g��!��z�V�;��Z���pM���:�ߵ�=��wl?u*jk��,Z��\� ���~ ＿�[��
K�'�C0���wPN������dz�E�(�DĊT����X@EDi"X��PĂ
b�*�
Jo3����|����ν�]�sm��Α�I�wv����>ť����W,��r�����*/���Uީ��~�zń���V9FЧB�n]Ąۯ'ϖ�t�6lN��G�	�� ���]�*���O�����U�ΘC$a'��eE��.c�՗2fToF��+��B^A+�|~\N��.<�ln�v +���H"α�U��O�y�/�}N�͹}̭���vݯ�V�!�дY{�el��=T]���'�d���xq�g|����{?*R|�l�d��}:S^�c�ԩ�޻�S{��Wg�=�	FG��gQYZNaQϺ�Z_@9��5k�)���钯x��w�qQ��7�:�|�Q=�eW��
'��07}ϐ�.f�Kv�����V,V=��ݝ	��ڛ+x��0�$��H<�^�yx�0�=�),P�!C���aݹꪻ���DF�p�|����,��1GsՐ3x�o�w�=<��#t�r,�����;������mg�wk���<7w%%6��U�u�8=*y�����$�L�Ï�Ƈ�����#���!�����6�$��~*��U���3{v�����[���x���c��V͒O�Ң����¦�����0�COJ���)� �h5���*�K�e[��Y�5Ap�\~�P[Ӑ����F�k�`�yjk2?�dH" �U2�l��0��U�_�V-5Z�o,��[-�lr
U�M4.͕)�RR������_�A� ]��tR9EL/#Z�m��Ub�T1��s�s�)��U2��v�H�E��c��q�r1��ט��I"e� �s	���u]"��	�R������k�F@��|��r{}��x��v�^̪�ߧw���,��{�r����l�e���u&��ꔕ�C��j�߬�9#o���M�qfA]�&��:�u:ǐ���n|�z5�+�d���Y�F�򒌆��j�y��I]:�媕|�ɗ*|�ew�FTVH�޽�Xh�o1Xc�#	v���r��L8T�Y���@u+W,c��K9��6mņ�~f�wkش�GRҿ��ѡcg�~�&�ρ�*#$��+���_�Ց�Ԟ]�ի�,|�5~���H�M6�D�
��=N9���[ɚ�k)�_�/����^̫��Qrn��_��̄q� v��s��t:���9�7G�=�ُ>I��"��*��4��ITWW�҂?n�Ms��ͷرs?������t�rC���ժ�.��f%���Zn��.�s���#�K�=�e���?�Ͽ��Y=���پ�OV��ȿ��I
�����X�hՁ�y����k�F�]�6�A|5�r�E}8���Ĺ���V��Յ�M6	�����J��kI�
dHf�^˦p�{@�{��鸒אI�͌��N&�yf�L �4����_^y��}��kp���dZ4[����.�^KvV!	iӎ�1�u���"iy7��T��h,�D��9J́����{9�����оݙ0�j~ڸ�v�EUU���EM��!-#%�	��Na:Y�A    IDAT~	�L��{� +�I	��x����x�E����rg��7������}5ǟ7��.]z�pV��Y�j)î���<y�Nvo�Fu���[��u�t��2r�gУ[W��Z�:��G�=a���?�"��xJBj�X=� ������<br�-1:3z��l	X�T�@�#m��@���c�/E�!�4�hEgL���,�VS�p�٢��u� �@5�Y�R��uX,�0Hw0�WU� ȂUQU�*��9X��q�$)Lf=�t�:o�?���h�����I*#����*���?���]7�p]*�7$/���$���IB���]89�*"�𩠷T�DŁ:r����dXu	�����&��n��&9�����Z�w���T{umm9�T�G*$�͂�f�R�e��Q�v��i^S�n�w�$�R=`&m��7H%���dZ�d�)�KAA)��X<��!
�Hiao.K�^�p5Gي��J�*c�P0N^Ns�8�,Uz)>%I:�u,I�l'�H�SŕZ�c����)5.���W���	���ܰ,4s���Lf4�D���2�v佔��
��E���dJ�@e��ibQ��(�jq�Ty82����i�h(��>�F��a�LZ���IH�.&���)ibc���qY��C�4R�ؾ��Z��Z����,Z�=�'�P�@�~WO�1:��9�� �c�o_����i����k4������Ϲj���q$C���}V't�y�<�����X�V^\�
���\p����<6&�YU��w�^$�Y;�",�՗d1��Ť#،.�Co6LD0��1�C��cևՕ�U�V���'�؜�U�dt5/BOɣQ,Au��H���h4�l�S��#6|ޠ�Ӫ��D\�V"q	X��~�(RA����ܪ�:�`Ѭ'��WZ��.����:��a��a�0��T�)�!f$�$�N��� 5i�V]Nf	lK��%�8I�a�0ԳX���"H_]�VNi��t�1��y;����G*��\Rnł,�
��%Hꢤ�Q���;����жm[v��S�U�Z3���#Q�'R,�$��cbW�����6����A1�6�I���@��aЋ�F�2vRqm�6YE��U�X�S����xF�+("	����R-��Wf�Y�=�փ��GO�%�,�)�01�#`$S��}�������O���%��1K���'�6���$-lduM�r�����v��HJpuUF�Si���J ���'�,+ז�n�43:�܉ X��+@cL�KJ/W����rW�f���!�R�{?�S_�U�*���pD��	��ۙ���>͂W>���X�l�F3�X0�͢I�]N����������������\���n���y��t>��:/y�n�PԆ��Ԫ�m͚5��݇l��l�[9.�JQ.��~�5�z�5���&py򨮬��]H"�P�AN��D�բzx�Y8��e��NJ9�XO�؜",N��2�͡-���9���Q����@(�Qgc��EG�ǩ��M:;ј��^�Ø�)Rqae\���h�h�+E�c��!f���T'�*:�b��7N$d���	�5��h�T}oTڏ^G`[*��m�Ř�b&����LY�:�J��k���9�Z��I��)�48U7��?�!�����jU�a�'�ʲ:�gjִ)����b�,6e���(x�T<�ͣG����8���Y0��㈦u�V��4�D�x:�ID��ш0O�qdS�O�V�ZD�:�͈�¨O�W}]��p��I'��������d9�FB��h��שq^umUՕ8�F��<TU��̚��B�^$��u=e�4��V�m+r2���PmB�*ɰ2 L(ѻ$�Jb��a����qg�	���:�]n������e������Iއ��͔��(�z*%[c��(��IK��'YK��T2F*Ġ�a6�U֤	�sj�&D�8�Y8-Nh�aL��~�lݲ���'�Y!8��tF^z�cf>�2��#1��F���lڸ���4������8���7w<��Q�ڙ��`4�rZ�u�k�t6	�K��{��oh�1t8�h��r�u��1��Y����nRf���َ1��|���*���̢���w���,Z4m��;�yx�0Z�H�յ\���#��n�*a�P�!������i[��#��؂��
������%tdgJ�Ƃ��ۻ�=��MZgT�'�ӮFU��jLf+f�d�ɪ�P��|��V<�"U��%�,�K*�KV�K�e1?y�\�O#9:U�ոr���a±0!�4*cP �%����r�&bD�!R2�H�HG�T9�nނ�r�6�%K?�s{��O�Y�l��M0RTU�+�%��?�ē-�֌�(��ĉ+$RP��5+_g�łޤ'	S�%7ˣ�o���e�)6�jwI�!ɔ|fБ�.�x�t4����
H���Rc2�N~N`3{���F���"c(�ӀA/N�4u5�|!Ud)ϟ��k7�"d��d��Iˌ�[W?����J}��L2��3���]餪x����9�3X�|�b_$+&�)�c2��xb{N�хW/䚫�婧���:�@�����aU6x}ڮ����vH���R�����.B`	�tX�	����#M���
�E��뫸��m[~Ŭ3�,�	����y��s-�9�@$�����_��c�RTr4FW�bh�@l��ɍ�����i�FM�g�=����ڬ��6��$�d-���f �ᤲ� �����[6�e�/��nZ4m��'OAn��d2ۜ|��'�\;��gN	u�&Gf��`UN��3�<��V~M] ���8�T.��Br��T��Y�b��)[�(�W�6m���({ۭ2�
x�ܹ�!�[�I5h��&.�{>m۶Q���|���l��̥�W�U�e����լZ��'Wn��0�t�֑5�6`йS���t�֙]���k���6{���tbX,꼵�kӜ��sX��Z5=F	8�?�x|�Z6��=-[5�w��f�a�PQQ���$��:�t�FUr��r�j����O=΁�t�։&M����SҺ�b��n׉ys擎��"�x���]�����_���ѦUN<�RK�JQ��Q-�KW����%�a��t�-Zs�9���Ԯl�m����G�=��J/t��Q�,U�c*�:��:+~��I]Ћ�j��
����d�\)7�ݭqٞ��-��pٻo��9���T�גJpf�"j�+� \/�e��MC�R&���fF��2�M&)X���V���_�_|N�N'�v�z�T��ej�(����;�H6n��O�ė�W�H���b�i�tL��u)��Y%�Y}��3�G*X���u+�*C�T����s����8��>�$�	J����1hz��Ia�&��9��6^~�s�1��-����B'}l���=�6n\;�M�'���t�VG~�X�~��2��=��%�X"??n�B(%77��;wa4�9�Us�=�(5�qe2z�]|��
K���c���v����!�>��|)���K����1c9�c��%�޾��O��ͣNg棟��o���7SY����"���E4L�V�<������8ruu�=�Y��N�ŀ~}9��#0�F gw�yu_z�ّ�^��'�zN1EEEEl����:���{2v�|��{�6iI�����w��g�7;7�><YŘL.a=��_�y�{2z��<>�y�{�aÆs���L��֮_�[o�c��-�����hކ��/��.ʍ7�@~A6�?�ʯv�ɒ�
����b���q�E�7�
.��&eɕQQ��mT���'�d���2�<^xn=߬���à!g�j�&n3���}���͘�47#�>n �6`��[���ʫ���>lڴ������c9�&����5[��mA(�'-ɷ�`����u�H"j4��m�U+wL�4R��9F4A����ḩFj��Ȉ��o��Gd���|��|��[5�g�Kӟd�J�d�L�LFd{H�ٱ�ѩ���`��c�*!!� �߄Vj)�i��	I���ܥ���D����ӪESd�Ԓ��V�#���Νe��UGZ�P�IF����&mt���Į�@� )�դ���d3驩(gȀs�j@/j+v�����P^������a����GQN3����ܭ;O6O>w��K?�	W~	F�K1��h ���)Rm�xk<�h4ء�gm��n�i0g�̱���9�s[.�u��Ӵ _���޵�����R�/�R�|r�[^Q���~��Y��Y�pd7�N,��<a5�*���7�k��ƛ�T�˼�35�e�nѴu�~�\t!U�Z��5��\uB}���ح�jQ2�Q�{=��䧍L�4�H$ũ����b?~��9������c�xv�{��߇��M��\�|�3}�9��n���m[r��;�g��=ŗ�~P.��l'S�@e��8���q6m�A^^b)��f�ʞ]��1m_p"�O}�A�e�;q���qS&_��>�������7v<�����#(n��ܹӘt�c,x�e����Is�T�Gf���e�m��񗭸��"�T)��f�c3h٬����
r���W^}��G�f��1�y���z��Aa~��������ګ=��I�f�>>�YO�ɜ9(�m������ŉ'���ƃ�M@F�&'v����R��N\[�0Y�l,~WV6��Ni��� ���:�X�!�o�Y�ɒ������&��hV�϶m�RX�O��_%N�t{�j����ih�΄�=�Q9��ߚ�I���/LNbk���6 �+H�� 㨒��!r�sٻw/�xD�W�lKl�jk�TV�),h��jS:�I1�M��40���E�����T��h����8�����9u<=s<�nUX��q�w�6m��H(D�VmIE��+���mh֪-{+�n0[S�&��@����^��Q��:���^m#��ӽ%������P�U��L,x�p�����pf���uTVV��/�1[Lj��&NM����f��vn?�Z���&��*�Dږ�1�ӄj�rͰK�n�9�8�AW����r͵c)��b�#'���۶a���|\z� J
�1���0�rT�S<YǾ}�0s�dB�x&ܮ|��K��Z�V#��*n��Z�_ދ�G��q��b�'�s筃�t�1<��B��!���J{v�HU�^z�ޕG�����5à��a�e}���~x���ɓ����W�Ե��19�å�l;;3a��xX�`/���J�=���{�h6o��q:���+Ը����9��c�={�|��,��-�ى?���˸��+:�7�.��5k���6�,n�|���{�2�[8��c��ڑD�q����?��*������/�g��M�W9�ڴh�m���d/fȕWq���8��2N�A�=�x�*�r�Q<�ح�;m�b�Z�mO<a �+�h�$�&'� �e��������*ݿ��}���Ha�XL��އx�̔W���Yiڬ����TD,��]�@�';Ksmi�ʱ�	�Т��N[�w�z���M4\�����e׈�I[�ѐ��1b��E��"$�j�8&�!��ʭ%}U�����I��q�ʍ��_-P6��gڶ�$<�v�Yu�I�km�6���N��PS���lYn'۷�"�Ӻy+v��&���{��+a��{X�q��fD�:����h �������xk<�h4Ё��m��eSw�V�Z5�uB�OY��8�\~g��F4Q�۶PSS��n��IsU��oY�a;���$R&"�͑L�t�H���N	�3䲾�tS��}	#o���������	�I%%/ŦN�d�CZC���i�!���&:��=;���8r('�J��z0l�m����B���å��3p��<1�	5.;��X�vW�ɕ��������8炁�޷�,��1Ƥ)c�z�6l؎�l���p:��x�(Ə�H�n]���)��_��� /��`8A($�m��`��s9�E��nO�}���<����E~���~ڢ�[aa6˗��ީwqJ�.<��$bI��.U/im�����ꡌ��Z���
*xI����!����e˸w��\p^U� �a�;�_}˻o|@��]<��Cdg{x��%t�Љ�G�f�W�ټ� ���3��@��I��g�Jꨪ*��Z3g�^}�[�;w^�q��"t֑�'��Ø$'&��q�F�aQ6|���UX,��̐rb0Y��ӄ"AT�aw8��������<苓�W��h��Mc9D�9elܪ�Iz��q-æ�>��ʁ�t(	%R��J#u���Z�����& I��8�b�����'$sǯ��v�tFu��&��X<�E�q��P��NO�щp�h@g��$\O��X�t:�R�^
�*	�mg�gӱS+�&	�Laҙ���Z���Q�K���j�6��,B���-R��^ֽ~w�z�O;���^o��O���]w���)��}����&e��F��E�hZ���zұ�q�=�F=�7��{|�?l!����5�@$A,U߇�t�z���e���*.���Ͻ��=��I�0↻ؾs/nw�PW��݃�.�A/���HH\Mr]˼y���5�~ϑmZ�ve��o��۟�&9���0aO�{��˗��)&iȦ����[�y~�T�~�M^^�:M[����@���p��ذ~+&�C�fMy��ix\f��#:O�0�鷙��K�}j]N*$��1w<�ʯWp����}�i,�t9M
��s�rrrؾ{�.n���&Q�����̸�f?�4_}��7�x�����'}��m����WQ��M�qˍC?f<�<-�������J`,���R�l}�e�i����_|�Y��j�1��{�hw��pb�.L�|=�.]�o�n������1]s�H��4�%�ܹ��z��3G������۟�WTB2eVvn!M�j��Y��_�N������t1����D2��E
Y�r\�~XD�"�L�H�����\Xr��+@d�iTϝ�i�����<���QTZ=���'��cr2N�޿�~넙�U�vR�v�����e,)��x\,ؚ5;��el�f�A��.X@{&(�!�Ҏ��H,�@���CR[A׮Gq�Y'c1ƈG�dg����nw�a��|��j���h/�d�!.�f�
����D؟^�ꝙ"���i��u�ɏ@#����A��;y��#Ik��I%'%&`$�I$�c�o��ҵ#F\˦�b�3ϩ����f$�&�7:��P,I"���J��hRm��ڸo�Dο�H���_��%��ͷ��x�X�*(�g��'�i�N��,)�
&�����m::w=�#�(������'7�ͻo}��3fq�7q�1~�c������x�z���޽�S����n`�̙;�#���q't��|+�ٝ��"��W3e��֭#/���6� ++����@M]-7���q:rL�#U�ޒ�@�佷f�޻_3e�4iR"+<>ٹ}�a*����Q�љ�J/���gX��*���"o,���l`���I�Ҹ�ݴ�p4v���9��O�}�ٳ��c:QVQ�'�E�_�ӧң[�����*��M�s1�%巆y�����{�:e>��^N=�$��7���~���}���c괛���y|��K�򪬬d�����ߕ#b��j����R�?�*���h�ɐ�Q��F�"F91��Á�ƾh�ue����j;2L�J�5��05䦕Vj�V�F�W���1/ٝ�v3�&��8�Ծ�ʂ�אJ(wWUE�z�bѳ8�������Wێ��k�YI�����djt�w=ճE�q'L�Q�\aƴ����R>��L:h�,O3�V�p������@�-�;�P4���v�bI�=H���}mr�z�w9a�E_G��/����v���w����b�dc$�
�3bLF1���&�F��¡N�F�]�$�-�6+ ���^���M�����&F�����t䦛����_8p��އ/V�B0�k��H̤;�a�ڵ�s߽x<.ƍG�'��M<�[WE:���������Wv�~S������R�>^�A]	���x����K���h��ɋ�Md�����mN����*iZ�͇�<���-e�/�����~�3���V��rA�^���S    IDAT�}3�����o�O�ݥ�.i���fL�k�\��f<~R���r<��9�����Q��g�]�βJ.�d �Nh��k&������������4oݜo%��̍׎�����GY��rv��C�N�(��e���x�i�ֳ��n��O������hp���rx�����1�6�t 4+#G^O����<y��\���bF�zK>YO��*N?�Z�2+�������)V6l�;_ ���PXɑI$�nBR�u�c�3#�e�XX-���8�t+e���byR)�%����q�h��ڨ萵;Z6n7�|g�C����ȑ ���)^u�lf�JJ6�IQ��ц�jS�)qdi�R}�e=`�"�':�Q �6B� �h��ܶ�
c�f5������I�b*�H2}�8۬b�7�7Z�J��,&���h�jg���6���{��ze�.�RV�H9a���G�uHI�NZR~E�(Z��
G�IR�B�f��nҺ2�IڄES	c�����V|��d�E,����ƙ�{ѵkg>��3�}�ZiSB�Z�_�We�<��|<�|����^���#ALF�j�.,�gŊ����E�����C5��S\܂ǟx�M��RW��D-�:O��r��)Gg�`�Y���*M�g�nlݺ���*.�ӗ�֮c�>��dc�I�q�������u?P��!�at����L�[�����`�Kid���;�ēW3z�Sfѭ�qd��P�����RW^���[�t�П�N�
��T��~ܴ�1�o��SE�y��d��P髢��%��0t�t�pg��X�H"�ř��`E5�-��=p8M���;���Ϟ8{�r��9K>^��e���ҺM:u�ľ}e����lڸ���B�BoQ�&�ȑhJ0�`
'�5�X�ą%�j�ƐdraDw�q*i��o�o�z�J�ڔD��_��2�A���o�mɌ�2�OFH|����M���@\N���R}ev3.���,��4_/^�tx�0[�X-6�Z:X8)����ɘՊ=\��Hh�C�1s4���!a�bqV����)�cr��6+�x<"8Ƥ
>C�
�4�t�:��C�#	�z����Ou����L�����!����;��QCa��93%B�*^
$%�6%�B&c�B�'�N$ɴ�2IU�T�j��rbW�$*7��4���WJ�6E��x"�41��O�b�Yp�s���t_�N��e�`�K̀B%QV��TS��b]���Y���A���&;�MJ%b18�؜��2"��P,����R�(�		�s8����'.#�HX�Tvi�$�r����� w@��zk1Xl8�n1y��f|�Z��͊��WZ��K�èY�B�*��ܕlW�����2�8�!�$)��X<�!��W[CQ�|Ճ��&T(��S��M��H����`���Bb�$�p��L]�h+
1��MF�$��D�O0R���� ��`Vy0�ܬ��FՎ�{�N��E[�%m+�MTH��l���V��f�
�hsdK('//��GyY6�C��G0��� I��Ża6�b(�Y���9�ƝylC@Ӱ�I5a5�w&���ʄ�_@���HT4%-�R\��1�����_̒%�R^V��  íע��jz��fH �8�bф~
�(Ц��l�P���I".ߓ�z^�^4D҃%ϭS�9O��O�Y,�1�D��P9NV�[	���@j��I�.�?��ڸ��h4�����x���a��c���\�k�(�xR�
6�/L�P�f�Q�%��<���5YD/��qO��a[]��H2���mBK�>F*'�ďV�AQ��P���|"��֘lЄ��y	��Ӣ%ɸU/4��mV"��GH��"���h8�N��*�LYjczb�89��� �D���\��K���b*�$�b��0Y��T����k�J�,�R��#�U��=Iu����������}�hն�*\$.u6jC	<Yv���,)"If��d(Aue�W��1��!i�ހZ<��,%�6�-�!u���<?���*���1Zͪ�i�A*�r_�8�T�o��.]����舘��q;��������Sl��ZF�a���b�z�UA��.j�X�f5Ҩ��aॗP^^FAA����T﷼������}2�~F��a%�G>��C� ���+��`�w,K}Ǔ<N�a�2?7��5H�FD��Z
�x���?�-���;��u�]���s�n�&�J�ƭ\�eٞ& ���T� �E鄴�����Ri����O+VR���w�l�i�<h�v�*�O�vB�-��g� �ĚW۶��'����G��4~@��G`���1��)Ŝ���F�n��^N�f5R�Z-�1:�N�V�E��r�Vm�FM��^�j&'YaA�9Y؊t�D<��a������bm,� �Y9Wd��~\]ዸX��=�<�ґ��Kᡈ�ejԐᰀ+՞��b�(�`&&��Fao�\�bS 'i��T�q����.A�,I}�xT,���E%��΢xBtiH&0�q�E���g ��Zu��h���Y�x�.l�,j�I��>�6�5�x9PY���P"��P���j�#f����`�9L8��b4+�L����9y�
ʨODբuv�l��;z�ғys_%�nJ���[�q��g2���

�PL�N�~�|�E��S��Tc�j�
e��K	c��e��&$�)s�M�X��-P
|�;�����y�ߙ�bf?��W�t=�E�I��[]S�Ҝ=.�V�Y�������T�X��s!��ld��$a)��b[�e4�1�� ��K���z�/�xa.c��&�-��j?w(�~��ly�RLF��3��S#����I7��;����w���o���ӦQ�u �=;,#��d؈D<ԕ�02�@�B�(U�^�N��1��G5�hD���� W�:q� ��6G6e��Mt�ԕ�6�F9Y�֗^J�daH&M�����Ț�@z���Rn�Y��������`8�EJq�5$�MK��p$�F.�������a�����nr�������x\Y|A|�H�a6��@F	bǶ[��$Z	����쯄�5mZ��nT��
G��Z�eڤ�Ք��ׁɁ^�.)6��ԸGz�ј2r_YeQ�Vg���� �#deۨ�*U#��L6JK����S�a�$�W"�C�
���@g�lJj���"�c1[`k���N��G���G�A �%+˭�]D����ς�������D\����A2��L�d�熋��`$���NC�Й�pՐ��ՈK*�l���P���T���kI�0/�E��\U�T{�XT e$�F����H��H��3# I �0{�pD�i94^Ф4j	�vR�8�tL����D�����p��,3��ݢX�T"�[
F�����Ջ'�������G�v���85���<��U^L+�04Ѹ�ɬ��]ѪUJB�4g�jdV�M��IM<� ����D.'ݪ���6��X�d	�ٗO?���8�v��n ����/�!'��4r�֩�,z�F��,g������詞��U�(�z�*��ę�'���Vj�~޺�UrM����	�g�e�M�.G�bٗ�+�-Ď wL�{o|DuE5g�}�Z(�����ƍY�r�Z��ԋh��нGO�?����b�R**��_�G��m�p��j�\YmM�l�yz.�vl������vBD�$�ϖ.c��u���pz�3�X��s���� ?n����.����篢��E��Nᜳ�*���w�g��+1�$�f,�<��֋�W�Ÿ��2:�?
V/�Q��ϪIs����݌��>��o�����j��R24�34����N���!7�� qxh���)1���]�4�*d�N��)�B�u2I����	�5���7Ʌ6F@i��R�NU�z*��PP>�J�Ѭ牔�~"���4����0a�~�eM�6g��],_����H/���i�ɑ7����TuB�����	�Ͱ5�DZ���z��x]Y��4F�^l��oMl�>�7ϓ����@#����_���G���w�����4�V��<m�/��"=�B�F�#Z9kW��$��P�r�	�0���2�HW��_hլ=vs�{����+���N|�b3��}�IX}h��)ʸI�`��x"Hn������q˭�Ӯm�S�'�.�E���������e�4��J����$#"�4K'��Ҽ��}|����i�>�Ysf�3r,�?���:��x����1�^�6g�s�`�'���{dg�0�~�67Gَ��H�����=�=�t���x�N:��֬^�I�[1k�h^X���%M�p��۸��+q��\v�i�=W�h�hY̅}��yL�0���Vs�Y�u�U�//e�W�ѧ���/k�oa����nN4dC'���HJ�dfi]Xi.��)Mr8�-?f���a��E��Z�3W�up�45d]2"�����W����Y6��:��?�ٗ�c����$�\r�xT��tIA?��O1e	�3�Fl��[�%�����$�gƥĳ�q��^��^�P����"_md�'m����O���$�0C�x�d�Ʋ����K'�R@�6����5-J����;���|�x���h4�������4b�6�HK�5���Ť^Gqp����9K���V��Ћ���P,�@&���m?QUQɎ��U��8�f>r�w��{���C���*�{�7iƯ�n��+��G�XG�)�M�f�q���?K��復R�ؒ�펣�	��q��|��X�)�X4�}�Jz�$�_?�$A�~��&��x�l'�p��{��������q�u7���敗g�M>�í,��?s?^z�W�|��>|�ϗ~�mcƣ3:��&??[�:LNN'V��yO�o��&����XLz&�>���b��7+'QeiW�]So����pB�c9�S�M8�`_�.�u=����9���S�3����tq��6=%*>�μ�`"��/�Ï�� �h��(&k�D2B2�u �-�
��-�3��?L(�
�G#��zFB�zv��HR͡$(��rX��l_�&�>�C�7Z��!}Ϳ-��C��>6(��W�E�ii���⃌���=��f�NU�S>�*?F�di 2��mҾ#�
2e��D�q���F�ng��վȗ#%Z+m�Kh�)�4#�V�=	s��G#X�Q�Ⱓ��lP����i<���G������?d�����.�.4��%�"!�^�2��yC=3�-�r](W��[$����&�R�,n`��"0�ߎ�X���ޚ÷�|ǑG���u?���s���q��WPPd��eK���x���4iR��z�:���YOp�y�qϽW��[��(��ͷ��0��L�s*�MY��J�>�lJ���Ȭxr�4j���v�,�6�p4�#�>LQ�G�1<j����ʤ�#�j�ilڲ�1��#H�����)��ζ�h�"��^З�%M9�j�,X@��c�ko�[�R-<�U�|�ݏ�{"�`�8���)�)Vz�_��a��r�'0���<u��V�����0rT.4�+���=zq��wPZV�;�L�c�቙��|�s��>��?�qw�R-�9�%����΂�Q�2t�HZ��L �\���Z�p��S5Zk�&S �FK�lL��њ����#Y95�j��Ȇc�tZ�\Ƈ�����N2�B�� ��U��p#��
 k��p?2��F��ǆ۱�<*:,I�)U�5�QQXƄ����0�4-Lf+�*�׋�.lNZ����-l����m���L�TD�%�)-L��$.�0�p8H��I��ح6[ �1c=�c�Z�l�b����'4jh�!��?��l4�w�o�_=.�����q͑�Yi,�h'{��C�HUq����f��LxZ�1-�U%�J�5E0���O>�O?��Qo�c�1��xy��|��+ο�4֯_��o~���b�ة���[\y�`�4�����n�l��@?�jw_���E�q�/<5g"'?ϻ�͝�'2``n�e
#�'N3�{1�r1�mX,r��Eti��*W��[�v<��(��Up�5��p������8ٵk�p������~nw;5� =��ۂ�)�	't�������%���s.&/[�A�|�n?&�ʠ��3~�ׅ�z�串�,z�]�|����С�������>��+��_z���|��Ga�mW0eƋ,Z�>mZ�@4"���Y��m֔�o��d̅��A�O�1��M&��E��d��ĝt���&�n3�F��`UF��LñM}(�� ����H��K2ې�Ҁ�*�j�����[���W���}���!s8�R,P�p���r ���b�Ɲy-"(RMRy �&a\D����NM4/,��9 �&9L�ę���ʡў�>!YR���A}e$���w�pXy��7*��jUD�EF��d��I���zh�Y4���������h�j��_t{�Z���1��m;)�Q��:���EN�ڢ��*�B�^�w����c#`'��fQ�n��;xj�#�������޻&���������k����߻��ѷ\�ț'�c�VN�ځ�S��㏾�Ď'�՗+y�������g�棏>b��݌{_~���F���ccޜٌ��Z��n��n�%,����I�	C�M.҉8n���n��%BI�<>w˾X�2`�y?STig�:+O6�θ�߶�ƌY�X�����t���l�RU�om9Ǵ?�y�g�n�~f�7�ъ���tS���s�2n�p���+֬��&�MY��*BA�*�7�2���/.�H���)�N�@���\3�f�����/����`�C���3iT7�F#��n��?�@"ͨ�w�Og�ά�@ď�"��@fkc��.�~�#��F�>���=�>�ZO��*h:��`�Põ6:�����w����il��_���05���<������ᮦ��#�&��J�e ��:md *w��,�\I���K�1�tR���D�ZI�v?��*���E�*�@��S��5�>�|��sL�S�Y�6���8K^���,��T�Eah�4�H �͢�}�xk<�h4Ё��m���w�b�bdĔJ�`8�EQ��j��+z��g����J��v)[�,��;#�\��b�J��铘u:�u�e[�6�N��3�.]N���V2���|��;lݺ��˜''s�����r� �O͘[��++��iۦ%^|����E��੹33�>֮۠��:�t�~k1�=|?z����=@,m��QXP�E��`�J�p���gL�v��s�@.4�[�������o���w������%�틕��z]��!�_����q��\r� L�"��#��0�_{������/��꠰�_D"g���{:��������G���Wʄ'7�����5�*��}
��p/����G�3��'	׆�{�=��~�6����d�./���'����d�Ky���4+n��V�6�D�I�#l�#.HI� 0򿨪_P��NӉ4d6�є�n{pԤ� ��P	ɹU�#�v�ܧ�X����0#F�B	�`H��_hh24E˙�m�49�N�S/�� ��E��"��$FI���U���M�a.�G�&�@������Z�d,RBBD�"��r�t�zT�˵�X'��ŉŃ�*/�F�YՌ[#�E14�[3�	��*+J/�n�0�L�g�44ѯN����k����u͟�����T��BSR�!���I����띪�@�״��n�{I�0?O�TUT��;s�Ò���W��!���K�p��iЋI����g��������ґL��!�s�\��~/���e���q饗2j� >�|5U匸�k7��[Fs���k�oV3h�eج0h�<p�$r�ѧ�����L�<�9��r��K	1��a��A���3w�{�u��L8a�C��ޫ�������ڱr�Ol�u�(ғg�]¬�sY��%:���㏾㻍[U�T׮y��9��T1�'	��,^�2Ƿ?Q����[�믽I�V�̞3�9Ϭ��S�ۄ�N�G��jn��
�_r�^�{��eO�V�v>�'gNeú�L�������U�*
 �    IDAT��ٽ� zL�p�lܸ�����*�`���+��x:L4^�C����z݌���� �tJ��W�F��c��_�z@s��|�έ��$�M=�~$���z+x��G[���� �������Ia���-��$�jT�$p0��p�MC�Of�%���*��3��U{��Ɍz��IFN�V�D�HK�)�^�[��Z��څM��n�[g��������Qӧ%bRT%Emu�DJ�h�
���V�&=&Tה���(�,O�0H)��Y��@"�|�ʝ���	���%�@#��K�M��<u�={k�f�x��HEu��q�C2.��6W!q1J6�A:��i�4�>�E�;R��ņ6���O���1�sU�A^~!e�p|�c��5���O)i֖�O�ʪU���)㬳OE��O>ZM~~!�vhN�S:QQY��/Q�޵uմj�L�BoڴI-��z�j��
���3ϡ�����z��2N?����x=f,%�
�>}:�Nu���az�>�x4��_lf����������b0�z��*`N��e���7M�9������N��x2��l樶6��}���|��]�����T�T˒٦X�	�x�Y�[��Q�������۶=6��c�i�OA���Wb��g�BHyO*��YӦ��(6���vG��ǟ70x�`��p���t�n�~��	I1]E�K�Cq� Ȃ�LhZ'2R�(7p��0���N����d4*�(c��G�xJs
iY*�_t3�agd,)��搮-�J�ʅ`P����N�L6L�y����}�d���2ld\d���K4(�&���~?eD�������R�	_]���J�R
�(@# �h��tHؠ���S��J��^�\��kvk5"�Ke�Ŋ�f����͈�bf��_}�@��=����e�������.��ϔ�����lI#@H�Y�J�� ��f  �����{oJUT@A6��IB����͝������]y������ᓭS�3{�3�9�9/���O܈�b��6�>�v��³��n��.�3}H�u�Έ� 4���g���u��h������8cԈt��^A�D�W�/8_�i�p�1�"[�aF)4��+���[l��- MyW-]-.�]�Q��������J,Ջ����N9vY��47�j�η:R�V���PA�]���f�jN������%1�eQ��=wUS�[,2�w"�T��Ř�SX�8�*C�aD�]�f��9y̘1#�E�*\�Ia�Tm	vd�7L�p�V/C{�
58F)�"�0���>m�U$�!�l�ŢL����6´S����>�샇|m�N	�dFU8��)�=R䪵�6�DQY��kנ�k�<ٯ\�믿>ꕪ  :'S�ə�K�
�b̢�5�O��P�i����
Ų(1��z����Lf5�g8����SK��64�oe
8q����P{b[jBhT��I*�1Mj���R�R!
|x�t�9��In�Y���b+��H�N��4*/iB��	���Cu��;;3RF����aT�$m�O��qZ>ä�*eN8!�V-&��D,2Yt�'�6��3N��{n�x�ď|��� �t�6����Vc������@HÒ�#8i�B��.����b	:h������4������Cm��ī�oxN[�sڈ��3�ZA��+1m:P���6L�u�X��
Gwa99�u\��ړ�����x�1yԡ8�����_�57ݎXz=hfBL�DC�T��)�y�HBl���*X���?��V/yBH��pJ��P��]G=�Fc�e�y�
�Q.�
r��A��(a'
��D��\�t@�Cf��:2/��P,�vC��؆U@���[S����&	��*�@ƶ�ȎI:y[[�T��^|�y�����Ï�R"CE��i��ͱZ8N]�mG��n@f	���}G�c�dz�t���K���O�:U�EZ10asji�	"Y�����뵇>v_���/_��OMֻL4��}���@���
ۙmdd���O�t�Jj��Y���ܛ�*щ��T��&(�e~,��m���q@3Y?�O	������c!9�K.�w�u� �_|	/��*\�0�CM:Q(�y���F�8�U@L.oJ��*�����ܢ�U+��sb��g�Q�P)U���k�F��.ݜN�����\qJ%��\�*b��?Dݍ�&�H�}@3��{���7|�i��
� ����4Ou�}O�oh�nͪK���C��"����Q���?�&��!�J!WX��f�p�Ջ02<�㏛�`��kGp��b��wÊ��8�c分@$���u������4��'�x"$L��a�@>����D�R���,׹�E�2E��[R�yy�w5��⨖FU�H�(J��l7�d����Cm�;R�3��Ph���EMN����VBa�/א+���كB�&--R����������B�D�Ʉq5ޞJf04�E��#�5M�tXN�S��7,d<g��p��O�x+V|$y[�G�u%0eKL@�`(Nv5�Є�
��u!��ݸܤ"��L�X��ٞ�E|��	@���	#=�bk�8U�� E��Tl��k��c2/\yIH�o�]��ؚR�.<�@H�O|y�~+j2kE%��@?���mIik�X+W�M�T@#����툂b��'&���r �Q �k��ٗ��MF)���������$����������۟ǝ�?�L�L�lG��9,ޛ�bƴ6��V�i����W`��{��p�	C���xk~}Ӽ���{Lk߭h��=�NV`�o/.֍�a�R,`xl��Ҹ�K�I��\�������G�?8?����&���7���wA��E\�߿�
}�e��O�,nL�.V���9A�f(�Z=�lnX(yZ'iaB4�Y�2���0b�Z�ZY�Jl�P7�Ne�5�6C����DD��!m�Q�XLMeK9�b��T4�D�B0É���4$�Vo��V)�teG� �^C��EL�ݓ�F��^%�f�8�~s�Qt-fBrG��?((-V��҉���>��UDC8��$�io�Q�)������B+���"�������u�%��T�?��֑���Q��D|Z&E!L�r�&'պ!c��[���kF`B����_���~�kD��m4��N��E_�g�L��0Ԫ��Q�ݔ�E�Q�r��-,�d0��;���o�Z��jh�rb[/{J�L��	�Ԍ ⱔ��v�j��5[mG�e��WF�~���F2M�K-������O9�O:]������:(HiЭ2��`��M�-�^���^�3Ͻ�T/���/���`�Sן���Z��
|J+�4������v�o-�����+E�Q��l�v��8�ĳ�f��Lz&�.Ǣ�����.�����{q��Gc�I�c��������q��?�-��6��U�,�w����^_�=w݃��X+����e�x��8��������~"O®�\�b���N;턟��gx��w0��������ٳ7����¡6�F��'������?�;o��h,��5��6��M����_��`N#��D�:�6\O ��ebippP
2s���
n��tfze�E
��C�(F`U+�~�/����C�?�?��etvL�rOO�?�x�Z�
<���bҤ��T�$�QF�mfy^'MCց��d�W�7X��2�R�
P���'r2;ܦ�?7&&����nl���'�Mn�H��x���*n�o�	a2�\�4�[�5"@!������&�
A������A�4|Ј��s�ˎ*?$��m�/��F�r&E.���?Vn�������:k� ٖ��r�0<Z�-��`���k"F&�G�g*ѯ��	���4@���U@*�O$�\�}w��/9���'�t�#�u2^����hvnc���7��e��8���`7È$ۡ9��"dXk��cA���o{c�7;���7� ����վg�3��8q4�zm?fNo��W���T��;�*�-5kW,���~��=.��Gx����n�H����`�]vƂ�����/~x���{�t��Ys�m�����h�w����!<��/�������{wv��+x뭥Xx�Y�����S�I+�q��>���-�`�p�[�u�_)�����@!L�1]t">\��r;��9\s�Cx���1�����o���*����eR��s�C�M1�?�ͷ��n<�=�g�~۽�a���׾�=�~�}l���Y��y�.�<$��	����I�C���5�p����s3���k�����{�ԩi��Oo�C7�Ϟx7�r��� ���P�Sw�TFZd�r��f�����Z�Ll��t�+�Q0(ڙ��1躁��ih8]
0L�3��P/q��D����M���7ax>0> �8�R<��}6D@���Q�` �RI@W,F�D	d	lhn�Y����P@=��c+�_?R��&#S*���	��F��aO�fK����/��-5���L�5��U���L�~/�0zx��GD\N��d2- �Lל��扉�	��(�Q����a�_\^�|6'��m��e?đm����~�.���Rii#���L��-�ע�#������1���P�utL���MF�4��}3���_���l�@�|6��g�(�;����b�3nRl[/����;�[��tG�t>�_6����X�G�N:n?�������k�쯟�)'��y��?���K��f�n���ݎ}��7�r%j����s��珽���/�t�x�w�w�B��Cq�e'��N�f�m���C^��������/�p���ŏc�9g`��#�N=���� 6�l|��#������_��_������q����������.�a����\���a	v�}7�<�$R����{1�`;N>�d��qɥ����o�;�7��{<�����F(@�ڥ8�{�Ʊ��2�y�I�����?Fh�iq���l�
�y�m��;�+O���<�G~�(�l�%r9`h��f3��h(��bT��а�p\KD�m�IL��f�:�9s����`p`������ՄE���ϠL04����`[�1�ՒQ:�64Yc�������r�Ր�a����?O�������4�u(b�p�%Z���k׮��'��C��+&��%�iԪ����ޞ��J�쉽S�f����hk��B�O4g�&q0v��S�@Mv�~Bd��`J�.�	%���D�B}�j���Hal<@���5��ţ1�̀�o�(�Vਃw�)��ϟz�^u�]���F��E��b�����K0�sp�9`,[F���/�܋���q�֫���
� ͧ���];��?��юP�����)#�������]��q���U9��qs���޻���z�*f_]v^��ۨ�s���k;g��
��U�z��e��9�.��������S���p?~�kq�?ƽw��֛�?x~�14�:8�8�{������~�8hG|爅b6��9{�'����8��SP�Pka�V/"԰f�
\���|�Y8�[� t��Q�������3��?�������Ǽ���w��s.A[��Rx���pQF_o~��kp�u��c?��{��T-�R��+�G*���?v]Ǎ�]�g��#�bl��` ���~l��F��Ǘ�W��k���ᒋo���l���As;�E�3ًD�(�sFȏgL���쇟?��:�(	�\�v �SD�ϕ�QbU��`��I��M-
�Ypy��y?�(`�㚒�1k��L�"v�&�|�E�~6#���y��`�������<���hK���y���G}�z(n��f|��Rd2�+f��*2Q{<���V�=ӆR!�c��.���E���C=""b��O�D ��UMir�6�ۮ���_<��j���{�cZ6�C`"�l�Q??-�cļi22X
�(��beWP-)��}Z��(��0�+����������Z����I�����굚����(6X�W_y�u��cx���8F��B�?n���w���m��k�yD�t�P͍vj�b�X.aZO�^���O��,B���$�W`��6�u����8Ds�?F��iHe���ޛ���8{���W�蛱)J�h�P�堹U\��B̙݉3O��W������]z���?��7�]�C��Ɵ�r���~8�ԫE�r�ѻ����������/�蘅=��'�r0��=p�B�A.?�=v���λ���*:;�bdd;��|~��?�K�Č���/A3jx����+�u�݁H�W�P	��\t�yȴ�`��E�D2���h�P��ۯǚ�+q��k��Ҫ:���`���8JgQ�Wp�����_Ǔ��9�G0s���_]��X�b]Z�	q��8-���|t�Ŕ�h-R�$>��#l���"6V"ՠ�N�p�k����Y�iF��E�8,��jaY&s�Dm��c
��!5V?���q�0��)+�_Z�T���:C�ai�ţ���}��c�����a��:���Z6l����}2?c�#�'"2�4{��;����$�{�=ԪlŠ��4%�� �g�|���A���O�w�g2)���X��-������K¾ҿ4�I#���j���^l9MU\o7tP��������|W^tv�~K��V瞿X�&5�L#�u6M,Ƕ�l�k�:�"p�ٗa��t��D�5�Ѵ
�/�wf��W�>3+�4��K��>�m�d�j�ۛ�
�;�/1kz
�]9�tsϺ/��]�L���a��Kp�¹��![�w�?��������?��%^}e5N?�2����c�`A��RE,�����Й���[���_�+��O=�Wy:�������^D�� �󝣰��O�ɝcN�ǟ�-��0:\�U`����w���z,*�&:2�X���g��c��#q��O�G�Doo֨����T,:|�<�쫈F�b�w�m�a��8����L��&
��E��s�����_BO�z������6ƭ�^����2��jK���(�8�S�]7ÑG-�'M��nD�P¹���p�X�uf��042�` "��[(���|@S)1eJ��hH8�D�H�F�cLL�X��&�{Tkɟ�af��ğf��F��x���>��m��N[�/��ii�x�Id�]����TkX�=�)!j]|@jG���\7�!X�y�)��� �rhDG|�(���G}K��="��H�Fܖ�ai�Ǘ�T;̋F��Q���[P�.~o�M6A6ϑ׌�K903�R�3��SC#L���;���F�}���{�:D���u71�v	�:�Py�x쉕����M&0��w8��ب�������/�h���g,3�L��"�م���yJ�g�]�u���h������6_2V��4����ȗʈ�l�}ݹ�`�0���r�[� m���.>�Xl2�G�NH�}y�j�,� k�sD�#D�ш�m��9^x�����pҼy8����~?���A4Ƿ�������X����C�x�bs�b��⋸�s������cOG!_F����y{����o�@[��o6sO����	y�1��ze��_��#�x�/� |�N�gq���	�	G]�r��`��OF4FsU�\굲�i�U`��MP�_�f�\�?{�G��~{�;���>\���}S;p�aI�<��s�jk���� �cU|nӭ�w�188 ��t;3�Z��H4.��������9vf��]��N�h�*���2U�*՚����
�/@DL���L���`��%��a�h2}o��x��b��P��oßP""����v5��;�J��V��2�c[���|љY�F��JzwyHjĻVE��C*����X$,��j�>�
�"�����j�ȶ���7������~����`�!�:4�{��`�v��/����
bѤ7����E�p��7	�m3��ks�kE ��-\qw#    IDAT����,�0���,ƕW<�G}s6��r�ǆ�'"Q���,|��*��G��ή^�	�5�8�Oa�o�8�5��y?�O=���O���f�E��҈���_L�j�R��������m����n03���`6�	ͪ!?��|ak��=�H��w/����YAG���@\�\���9��[���<�*^����QG��ޡ�|��/�{��8�����.������1'��7�|<�^��x�gpɥg��7�b�e׉�
�h<�8i��p�9��o}�}�x����pŕ�a��Y(l�����|�E�r�)8��k1mz��m\y�O���^�'m�=� Y�N9mF��8��s��Wg�����t����Q�d�$�0g�4\��{����7���?o��=\p��������30��� -�6�o��!�-_�D*�J5'�X�"C$�iI8'X���E8���W�Y0Y�)����Z�ݽ2�M��vF���[ ���M[Q�u02�#��]��c �t��C�-���M�p{du�nF�q��T��V�"mB�=��h@p!F����C �����Qo9�8�X�x��yTK��υ9��e��x
�t�]����8-��T
����bUT�oG���k��k���Lcc#�3�n������ �d���K⶧�@��H���(!�,f��@�W��P(��]�,���10PC8��լ#E�7�O�u�UG0s��0,_��H�y�Hd2
������^��o���:���h����i���(�4�R�\�J�F�*t�O���2�ʰCI���#�@2u�lm�4"Ic�A�8֪�R i�5sF:� ̙=���y<��/�E@�M6�G���Q��o��_��
�n�XG�l��F����{��1t-�D�n}S{$ �G�U���݉=v�	��|V�Z���pA\u�5�5x��q�����#x��O�^�l&�Ai��~_G$�����ǰ��������y��b�-�����һ�ʫo��cʵ:����L��ep�1�b�����?��;n�_Z@�\{�����:z�f"�o��X�j�0t fR�*����!�`W�Bᐊ��8xϰM�'~23,ξ���@P,�^O��34�r�YdY��?�]�E�\����s2bݰ�]��p���8�W����bjvS��~m4[�x��F�#tW��y�N��ԪS�~��h2d��F�j	V����pě���8���h�3'\O�+FZX��G���E�@b�[�4�(�q	�b�`� ��6��)���J?
��\�0F�FA��g_�r<tLV@'���Z�F0�9��E����D�aZ�snk�B�X�� �J�7����w���i�����Zl�cwfѢ�c�ol'۶�aǶ��m۶m۶m۷���|���5F���jα��\��6���U��S[i%8�[�߶����ZKO� NЉr��X ��<�� Q2lh=''�F�`� �p3�Mlsc	5zv#��_}��J�������B�hOr ~���W�����"��ׁr���h�C�f����ΐɆy*���P�o,��~����rr�i�&�y�ݟ^2iL����	`ɴ^{��$}��`�ؓ��`5Jg ���ȋ�~F��2������Ѓ���bQ��h2�B��\ha�p,	�@k:��V��.��QZ5?���{G~�yו�-׉#�\,�_��X�nk���5'>BYh�'�vK��P�vc��E���ݸ-<=3&�|��c�8�!}S{#v`Xb�Cݕ�-,���d�2N��+S��c�ŉQ���Ё�OǉR}��j��у�1SL������B����2kE2"��pC����d���A�}3�-u*�D��^^�&�o��(i��*P����Ydz��-.U5�h [��%�1,��m��9������CWD:��g3��]��5BL�HJ7����b���Ę���1B�۞�.v�
�"�a<�a�d/��)hj��R����W�B���0�ٔ�i�eW��Y�K�6�R?�J�~�� LtW��V�"C]@���Y{Oa��/I�j�3X_�
,.������:�C�y�f�5�鿊��)�7g#�,������I�?C���0���J�ǉje�$F�z_���aq)0c%6ܙ� F���svN�BW���%�k�R�џ��O^ua�bK����s�.���ZM����}�gs{!�N�,c�V�� �Ob��sT{%�aѩyF���s�ĮT�bD
T�I7�]\�e8����a" \�N6���CE�M�085[��A�Vr��u$U ��,V�!"�24��{�*��K��W<���R�0Q� ~�H#_��Ʃ��F+��2qQ��i��������@���jj�
 L0nuyi�ʠ�B#�7,�+�Q�$��Po*F�c�-j��Iε�W錄?Z�T��oz,�07ҵ�2-�`��!_�\�Uh���PD>f@�=ĎIH�k!�1�R�}bP"�@F�-.ɗh��ex�Ȑ��CaK^�ը����n��2̥���yڟYa���-������W�ɾ�Q�OՆY6�|�l�WrsQ%6ZT8�&4��l�&�)27::��49��k�<Wox�L�}#���ghV�O&#�Ȧ��6�O�Tv��.�-3�N+�{.]�����M����^r�*~WH��S>"�>Nbt�����p�o��xRc�j	���%�1>7b�~�f�Rg"ԥ�r,�G�46g��7&�J� �b�p���bjM�FT��ק�����7��ч�4������v�r�r0[�T%o��{��`ޜ�j�!4�`�$�T��3�I<�uI�<8�t�H�4ޡRU~�6h�#2.o�4��Թ��d5�AƾL]�E�;�:*���S�޲��M����{���(���^���$�����1a�rf���m�Em�Џr�i����� ޯ�ش��/kb�ٛ��V�sRՂS�(οtd*���T]d��k�E=x x������"���)H[p=Ё�#���W_���q2���r�-eRi;9�ł��J�D����R��B�
9\��eUI�p��X��%EN#��B;��������L�� �z��9�(آ���C�*��_�;	�y��U,�<@�6S*���"���:j?Z=�9,1>l���?�=�=�2�+���4~�U,{�� K��[��3t���#Ÿs�N��^�P�qE�M�g�DR ��h�/�v�ϡJ���h-�U�j6>y2�膒5{"��[M�E��� ��RR�CFE��p(T�����|����ۼ�	ı��N�7	7���o^�F��?	?3ڊ�l�6f3��!I��3h��I��S+�OA�x���r�zZ��YyF�F %	%�Ͽ:��U$X+�:��w�v�\�'�Q` �`��`��ը�eӢ'n�Ϥ���Eın�V�G�/�_H�\�2�7-'j��{��;���@�}��4�&�Q�7�����^g�=��j��ֲ_��C��|�V�(�j�7A��:�z����� 1HdX��U#�[�Q�b��]����6"2WeX�I��:+�s��ס����i�[k���ڷ���5k�I�_ā�(�`&r�d��'+ۘ�ë�����$��g�s&(E��q��ʺ8�*lJ��^��M������^�0<+_.#h�:�X�_�2�5�ъ8!W�c*�2�7B�A/6�>��*��P�#��O5��S������6P�D'�XZ9ډ8���wi���Tg���h�o��V�#P��Z�!؈k~>^bPd���E`�$cI@��I
�z�v�Z"Vf���4�|h�uwvv�#ӷ�<�Mؒ+�}A8X�s�+
���ɴ���ڪ���6 ���Ȣ����-�(Vqd�.r���E�G���ȏ羶�<k��7~.r�fW��"��_��b�Kq}7�x�;X�O,���R7h�]�)�C�Z�>�XW퐿�O²vu'��eϡp��!�>9E��y�������!2���??�r`s%��R�㠥&�����F��3��_�	����$�(�(���z˼�'�H�T�X@��]�g�����y����R*�^�&\�f�����̍� �+�p�77�5�ͱ�^g?���e˄��Z12�'^��=Hi�ǂ���c`j@����t\��f�����9���r�N2��#B�rs��K�iNRMe0A�g�ZZP�ֵ�f�c����G�?�mՇaVe�K�4[㳓W!%\ԂQE�/�E|A���i�����y�  �:��uv�͒ EY�ͦWP�9P-�bݽ�^����Qw����W�%Ȧۂ��n_�~�q-lj�j�9Z#�`�D�B7>�����������D*I`IR����fQ@�w��T
�B��`��R�D0:�F'4�V�o���2<l�����Sf�A���a\S�D~C|�L@;�|�?c�v�N����%�����p �.��,'��!��l��7E_��g�:NH�f�x]ʨ|K)�(,��@MB|��r�@C}ҍ~�/Y��j|8xxõ���F׿��Fh����0�K�Exb��Uj��	ssn;�Ɗ��F����}��͠��bn�6�@Wz��R,`�ͭ08&�p������^8����k �0���S���r�5u?��D �?C�I������Pq�	�n��k��S���z8�d�c�˧�X�'+�v�\6�m{���&��>��j�I4�@VJ5��������(3���:-O�eH'XJ?P#�g{{�;�EI��UaBc���R*��Jl͛2��2��q���8�w�v�Z�d��ŕ(^��*0�+�RJ|Y9����庉0����hPj�5��=f�V�@��W\uL�3��]�25�*�o���j����R�u33ꮥ�'ræ�b�`��w�i2Tx�G��i�)ĉ�2�@A���gjA_��N���4p���H�<9PDT/ ������MJ��C0 ��Z��	��?�V�=�u�'���שZ�V�RO�.?6%Ⱥ�Jv@��.܌��s؂-������1g��a������ �V�n-=f� �K �����jL�9�j[�&�?�l5��F��dm��7!n����	y�)Nv�ǉ��
}��44������������8��EE��ة�X)�CW,kEƕ^�<�\E:^�(r�)��C�����H]�5�*�=$���sh,?ӌ0�a[VƠ]����؍��P��|}p0�%u��� ��t7G�Q�ךU�y+��A���#�a,�����G,��C�ϫ��$)C'J
K#�5��ye��sMx���H�a�f؅V'r��{t��
7�# ���:{�W_F�f'�G�0Y��o�0̗��"C�2���A���,�Yaa����\K�I~W�6q�l�K#�;�1�Y�G@=S��7�^oz�'��~B7�tM�_���W7]���Z��?����}R���-�G-Y���ۓ�-Q��"pE_�6�3�7?�@��C���cy�?���+K%���Q�6z�I1�X5�&�/��L�iX�b����:@Y��p���zI�_�ŢX-�2��"mʞuOX��0�S(���k�ɤQ�I�s�*�����-���ם83��`���r_v�b�t�`re9���qK2v�X*6`'�km}��A- �7�zCwNH�O���D���i��#9���!��6U'7K�J p8=DqB$a�$��Q��a!T2�jyS�v�^�����!�	u�_�1[���qKs��6{� �huÏ_ӡ�g;�F�Q'�k��))�q��g9�n���0F0�=ڔ��<�a�����g%�'�iaY�y����#�VQ%]Y���]A���c��g,��`Z^4�Y,�̌-���][����ޗ�3�yJ`�d���Lkt����W���5�¾0o����jFhμ�ă/Ah��3��ً����œU���A����θi��~�@��A%�m���\��)�0f��@���b�:�m 9k���}�����U����?tG}����t<���6CX~fN�-�$2��%�-�7�VG$\<�I�Qs�:Oz��U��%�x�" P���,%��GTW�T5��`���6��5IA��1����gYX&iP{s�G3dS#�ޙ�g�[S!�"@Ê�`������]��ݸ��Q3I6ۓ:�n��Bӓ�櫩Q̓1��lA��5 �5���[��Y�ˁ�l�+c�����̅"gWhR�h)ը���_a�s�(Y��2�0�ܮ�ېͪE&��g�κA8w�r�ӭ�1I���U�fƆ� ��T���B�?�,����Z���1��Lk��4'�����i��؍Ϳ�Z�,���#�F��(�M�R�&���ˁգ��Uj���֩6�֩��㶞$��!�����FH����F5��^�E�=�ם|���.VR�"��l�A�@��-a���W��'�V'�',�i�z<v���b:-���}����m2�T�o�tn��^l��+ӨX
TWYa�� �� *c��e_��Kx�u�����}�����`���$���Ȟ7|�3���[��u��_xI�����l�0��nF��y@�?���4���0��
���@�u�o��$�{����С�'�5�����Ֆ��R�5 �y{��$9��1�f��bv��e�X��C����j�WXYXȁ#���e��̜��$TF����Dݫ��}Q �71���?xɑ��U���	fU����������� D��UB\p��9,z���Z3D�p����ܡ/Wi�\��aފ�C;c�X��I��Nŭ�=���Z+�3�Ϟ�y���iYumq��_H�@���j�/ҨJ�0Jv�i�6��&a���vtBh�.?��2�wSj3[XC���֩J�#
;r����kpB�Ϳ��ϩ����AA��BW�`�����eʰr�����l֩9B�Yk=)'Ƚ�F�-'0�d,�5g�/664sb�at�mC�~��L������4�{z)��h�[yW!����c~��B\�X���z7ZQ�d�%5mdTRQ��s�r���#h��G,p_Q8�|����g��ieT�+ �.5��hd!����2E���m8���_�mi}.V�2
yHmڣ�l��o���Vh��b�B�u���X3�=8+sFcd�L�Y&9�e�A?�ʦ�Ȗ��}���|��>�zڌ�>\8�@�Z�8aH�����B���GI�+V��K;D~��Ԯ�q���4�^q�Ș�(iX��8��4��]ܢ;E�	��;�r�t����\<�Bp�uq��P�20�|&|N��y ��2c�x��n���8��43���z�P���ȟr[�Q��@��k
�ߤ��Z�6vH��=�8��{uK	����/�?���zȟ**�U�ih���)��[I���7z�����7^/��d/�ڠ��%�q=1{Q�LFN�U�"3��(U:��X?̬�Ns�1��W���5/��w�Gpd~�Yu�Qg(d5?��ϳ7Kń"�~ ����Eu��=X�u{������'ht��М>�6ˠ8e�@b���i���gr}��j� ��j��������e�-�� ��ܵ($�'e�Dq��F8G��}�ͨHWw:��M_���64�/RgB&��Ce��������6@��6d��N�v!��=�u+����N�6�*9�ԯ�z	L�����ӲjS�����0b"ç�O�)ň��ST��,?al������U/}�j�?�ЪI*�E����e�x�9��ǚ�y�lZ��v�vr��Mg� 4��(T�C��x�
����ѱ��<�}�Fr��"i���'��l�2��n�S��Ny�}]+G����e�/GAk�gUXP�ꑌ�Q�l�AQ�f�ID:�-L��EmGo�ϡi�z�3�o�GRS�}}B�(��� ��1�{�*��L2���G�ܷ�i=	����N5���jb���J�^����Ҥ|2F��3�N��S4�R�x!	<e�( �F�cdVJӛ�ȼ�&D���b�����ty�Q�ρ�?d���8^��<O��^�$�0�{�ٚe��?��C��epc!��)������_��˝����L󥷤d��}����ȏV�"��� 4x���!����L�Nl؆2����Znv{m��+j�]���Z�~*/T� �oJ��X#�T�� ��ȱ��Ug�vpȟ�,��DU���"�J'���#@�r�X����T�b!I�:#k�x���92,h�J��P���]4��A�~��� �R3B�P�%��hc���y�2<�D�h�L[����G�h�h8��R����0#r�q ����9�%����Sࠦ�cidC�o�x��$;x�ǽg*(�����\��-�7R:�G�����cgЀ5l,0j��85�:$w7Ъ|�1�:k��]|��\h�0��^d@��K=��Rm�����A4L
��l�{1�'�{]��{�<�����sXsh�Z2�u?3s⫟�Ӧ��r�tf�%��M����2���D){�h��6l�������1\5���v�I��d��n������{::�՞�N�5�c��C��u���D�&u�r-���6iG	a6��d����g�-SU��J�@D�[M����Ây�<7�2�p�Z�b��ذ��;[�iY:[?�dW�Y}hВ`��X\5��&�Bf�w��7��5@q0�Mj��L�Al����/��\+�q�_0����S)�-l9��+��q�&��A\� ܶXp����7����('u
�h��K�hڇ�n�����9�L���x;�~�R��2r.��(��o��S*�;Z�q�Tv��G^�0�*b�`�-�p@AX
"�?9`*��1�~7�d�bɃ�r�~�����HvR�W�������H�V9qJ�L5Z�Ժ�Z�J�I��N�!�1ɑ�}.օ���'b�ɮ��]"~4��u�����(���Z_D��ja��1L�	�,)\��C�<F�|6=�����*c2H7Gk4kaZ]�
p$"A��55;�?�w,3��4��/�gc��G�b`f Y��]���@����+� ����)�Br��k�_$o�[����(ε0�;��ƞ-@\_��Ī��y��_7���h|�W|��(��s���O�O1Q�����-�2!�&����p�U/j�7z�z�&!�����Τ p~����N��DK��K�W��DruEL���t�Z���`-L��o2��:)�K�.ç�HXYY��D�Ɖ1���m{o��1�+�A�Xe�����쥓`��)S�)1��*�k��ܘ�0�97,�/0��
�a�(�n{}��,�>�Vy�@��nE��S'��db~: ��`��,��¾*��u�s+��uɕ7𙙺�fb�me���V��Ip����=�b�
%"�1���Rͼ��<��2���,m�J��sv6�̖֝��L%�*m�O��A(�q+�s@� �$�c'|La�����o����ff|����V!���Fl���$�6o�S摃/a,Д�	�QX��"[T��]v�Y���]����U�9*Z��3���{��2��Wj���k�����*(�v����V+ZY%NjҎ�c���}9ޖ�u����F�?3ns��M�I���3���
�İ?C#�U �#k_D�Cp�Fŉa�3#�#+�V1��k�|P*��[��	D�4��Qi `P7��0�^��Dmߠ�S=�����&R�FrJ�ܐUg���
�u�ISL��)F��]5x�^�6<g�� ��*�S�̼�=ۗ{j/�W�f��2;�U�B���'���,��Y�2�ɼ�jwӺ<�#��k�RFǚ�{���=����Y�ӓ
QV��eʮ�;qPS���k5`w�V�]C�J�(2[#��HH1�MJy:?�5+���� �>]��D����ѐ���D��K��$	�f,5ID����en����,�����a�l���|YRbH�]�����E�����C��N.��$ ���u]�����F;؃5�<��Ƣ��؉��Y�ӷw�2k&������Rﱘ��;g��H$��]c��x�O)�]���uI"���@45�s�"�$z�(Wf�-��)C�E4�G6}ê�.��V�`�v����r���:���D�^w� /�2On�x-k��;�MV.*@k��u����`��)�J������_JY�)N�n0Ђ	��Av���.	&_Zo#t=<�O���țz\7�4�M�F��K�X��^f�&D��;jb7lN����#V]����Gi$5�1k�!�C@ Ɵ�˖��U��L���Ƨb)����ً��e9jP���¯�/Ξ�X��>��)"�*��Ɯz	��N��|�w���?e-����70R��hiM��=*R�>�8�·��y�T'Fٝ�H*?M�����gB'#���lz����l5�,�û��j"^X.�*],�h,Zz�y K1gz�tQ��1�R��SӲ�s���Ѳjn:4��jA��=0Oc� ��}��2H k�{[��F���b�F^��owo/|��Z�@�$S�j	��r��O�����~�����H-V����{�Y�����Űw�HLtc���-V��E��Z�stn5�b���;�i!��n��t%�'�u�|Q���0�7���ܭE3k��pi �`���ild��F��ٌP����Y��ZK2��3�(��� Yd�s1�FNG��l{�a_#q�M�����.��2!��}�Gb�r��������w�A�	#��x3�N+
 �B3�_���*�(8�\y���=��;1%���s:����Q��`��Sa,C4Qvh.sB�L�[���i9�z�gQ�����.KRC0:(�������ѩݐ�hW��P�J����YW2���+#l:M������l��e�T���	3��>���}N���;*G9H���3j�d���4#���Y���+�h����c����&�L�	�:T9��g��Xq�2c3ȯ���F	��5h_�}p%U����m�_PC��g�����a#-&W0�+V3�"�S�bb�Q�x4�����V�Q*r��x9��ݺSF;��)sJj�pWWț�+E���G�
���w��wϷK���F�W��`Ԁ7���`3��r��t�L)��I�~�.��Ϸrr�:a�<����/(�/#��#C�¥K<��B��ZX"�8L���eHZRT��1��vv�����D���Ud��Ԟ�,�6�����I���온��.�".�Zڑ�LФ�6&���MN�W("1f��hs���[R�V" �m�u�W�E�m 	��/�bi,bHŪ(��#J���&��L��CB��4,��P^�G��2_0�;ӟ��T�;�q<݅Q�sG��oI�B9�..jW�Ųݦ��nEv���&��۝j���N!��@e��7^@@^1�|���*1ʖl�q��+��e�X�p��Q�~�P�50H���.�ǤX:2h�9G��Q�U	�Uy�K4;����E<0�ÎL�v1T&�3�ږ#� ��ҀSzP�WJg�\3d��0R�8��%mϒ� 
�i(� cN�d����Ō��.b2�P�����~��� i� ���g��e�V���Q�ع���I���~^~�~^�i��MOڬ�����4��O���o�댫�J܆��������}b��4e�`>�c/q�2�#0��-Pr屆�@?-�v|��7��._ԓ?�y{�"$���=N� ��AR �cH}k�Q%ڤ����ŧA�y@�+��pq��5��1#4��7�?�P|`�B����X�3+!���t/"�ӿ���J�nͻG��4�0��!����S�ʴy���u�y��2�6����0�Ac���j��N�M��HK��°#q��D�͊��{�T��}pˆ���k2XP#�=J�'�5ˋ��"�e��kb�d�`ԋ�H��yH�&
���V���uǍ�ò"���O+a5Wm�?�o�7lLc~0��r���v�������ގ3��~�4o\��T����h��L��+��[��<��P�M�p��F��x���>�M�A[��^7s/.8vQMB��FG��E��ՠ1�nC�" �Mw��W!����4�S��6!4q/̗���p*�D�J���j��BlGe$��L"��:<U�D������Uk�7S9`T��������T�&�ݝ7��˙��cs�Ǳi��_�V��$��d�o����$/��,N�\p�"s��1�k[��������y���	]��/�R%007��̈���,ae}g(W�x  ��I'D)+��^~�d��etMeb�?�6�e�� �<2�𸬣@x=����$�i�k�N�^���0��qW�'�^�������V�#��K�k�we���ȴYU�؎�	�7�:j	��O��I.��]<��ٯ(�ю$��nH��<A����ʵY�ZX�DQ`���Uֱ��F�� 1�m',IT8H�BHz�X��d�_�'+�9	(�!T�1,Q�j�+��GP�<�W�&��ڸ*$<��R@��8l8�ס2M옑�p]i�
塈� 4NcQ�*�d��B/Dz�]�f�r�ht�������A]+�A|^^s*x$�zJ�t�%�X0��i2J��^�R� �GJ���O�:6����m�.$jL�<�:�M�Ɉ��PA� �Py�1�J8�U��M���b�O�D=�/AM*BjdD�o%F�`��_�����K�y�Ht��l�E;�gb�i�YU����셛�,H��9w�#'�B����?�.Z.E+-(E7��
�i���ޯ+��t0��ű���|�Fg�� pЏ��*Q(�E1�,ҾY��K,���Y��$ڄ�pR�d[P���7��U��	��sDJm�Ȇτ#�m ����I'�n�Z�`!�J�h z^�&(<dW� oj;a�U�V�X\���fa���^`���",�#H�Ѝ��ج¬݌Y*�lk��4�Yv��W_�l :��8�E���ok��&��m��O�m}����%ѿ�� c�8$��7QhP���R��#��� �W��C~�$����Y��,�"�Q�۠��^�!�=���ĥ���vJ t@C�R6Q
e�l6,��I�5� Ӵ$��C��HH	f]P�٥�Hoo�[���)���>r?���o)_P�OxpJ�U��`�f+,!�$�,��\%zX;G�!����;�� ���S����I�����Y�U&��>��vUU��)61���Q��#�O�+/�D�����Hޅ)�pd���]4VvE�(�R�!�1�988x&� � x��Hf>`�TP>Tfkv���}�u��g�,x3��� �&�˲.7�OGUw�l��fc���|�XN\Ü��̑a�xt�S�	7���&��ݳØ�'L��ܨ'i�(�4)��-ʑ4�N�6y؁�i�:idO��n+���<����K��V�L�j�̸���)Nr��q`e��diiI菉i��������h�V���	�m���m�1p��;��g1_���`^����:�y��ɹLD|.v�ę;ƥ�F���O�(h�f��L�4��Dy�z$m��9a�#���4�y�|�ȿ��I��f��|���>�r�?D�3OL�4����p��$��X
��IF���Tu7���HG����`$�,�II��G�
?���歉s�p�����00b�}�Ǚ�����V��З��������%�D��JGEʖ;͏2�<�|���z�J{�@�F�Z$��=;O4�g��3@��mM��g����_�ѷ�9�wȆW0�
��Ck<�Hw������ Ω� �����o-*J*�6��9�Z�(���-�g�o<W���T_շ�ō��YEw��Vm�!���}E<��6[s�v��Do��D
���^��a���܍ß~��c_��L]O�k�k�����|�/�/��;jώ+�1w��G�·km���֧f�:�+�M�-@��Ϥ�%�;3~f�V��y�`�;��="����+�lou���Z�Z�7�Mv���o��l/ �n��E�wfO�#��%�Oo���<J<��7Y2��Z�'3~;"^�#�S�h���]��BT���7a���3�ɴ�F�����U����:�z�7��͙���\��������$A���6�[���QR�ݡ���O+pǋ��̡����\ �ԈT�c����!=#Ԥ���X^ZiU���|)CT�����z���#��Fl�O C�bР����������~����P����q��O
篷��ÅМh��Bj'r��$	�2�GE4c�]�I��ⷕ�x����v�3�?#σ��߸:.���4�0�����?�H@�HĻ���gg{c�nþ`�$����4��X�	m�f���P���
\�ŵ.�`r���Ķ��rEV�Cr�}��
Ze�E��ƣ�S��҅����o����w�9H�O?6�M��d@���5��<��H}����UF� ��v��R�r�EB#��Ɗ��^�D�7�u�6@�:�����q�xV�?��}?:����i�w����[��}���[�fzΫ�`��}�!�i{��I�D���\�<���?��c�*ͨ�i�v�vr����Q&�I��l:�ʅ�8���E]gp���y $��+�A?t�����]ݲ�Y�},��=ZS봆��<u�v7� ߯�ϊ�s�Ϸ�J��������s]�j9��rM���'ʔU=�`?4��y:R�7��y�Ҿ�h��볠�~dQ����x��Ie����?��n4o��.���0�S+t��8��wLZ�g�J��x����f�~�8Fn�S�������/yme�7��!;l�MHU��v+n�Z����kb�#d�>�\�V�[�W�/6�nW��g����݌�F�Oܥ.H�{�?�W����N�IM�� &8��$�,7��a��#N)�E�"eI��� �,��՛���,�ٛχZ�	��[���R��`vE�9B���T���ei{���T:�i�L>TQ.Ѫ���w\�g�b^d"LoG���Kn$�O�iH��iA�0�uD��=#��Y�Ir��q��K�H����ԽUW�#L\���������,��C���]�gƓ�B�K.�L�2����*˦a����GB��2��.GX�a)̤*����F�v��=.n� >C�6.�8�W���_�7�p)Z��9�l?e��5)�;=���=�^s���!bQ	���&�����W��!k��'9�	>h��I0c ��R9?Q���\�t�.�3�ZW#������$��:4]�z�j�3���X���T�`��k����Tr��R��t��1OX��f�A͛TM�3ytV�hD��I6�L���#wZ�Z�ANH,���u��E��CT��}eM=��*����H���:��ɪ"G���n |���Y$�3�����&�\��Rߛ�V�*�Cvj$�� �5���݈s/��do���x�����������b�m?,�m�Q���c��b$�Ӑ�k��0W�>�������ᭀ��h�����@T��̝�������$Jz�e�	SlU� pXq���"��C�SM���[m|��k���9P��HI�d��X�����������X�M�í������8����n"p��i�6�n���u%|&�FA&:PAh�S�����}�A�{}3���Y0���p�ڄ��\vޯ$;R&�$CP@��H�#g����4��g��Hy�W��$[�B�m96נ�ޥ����i�jJ�[�wm�'Em�D��߿���v��T����-*����!uʅUvgѠ��C4�)R�S�"�s��	f_�݉����MD��@��b�߽Sy$p9�=�UR���drB���X��
 ��[�vT�R��Q���[s�f܁�΄�W��հ'X2�5��ɦ��vj̊�5�*�:����,q��� �~�����j5?2S�Cx(�		!ȄO�i��l�<ѵC������b��41鄅[A!ᶯ��?A�[�Pčɷ�6�߻ e��By�&S�x���ܶ]�5�;�3<����}��6�Cw��G�,���u6[������B���AW���n)	�v� ��ھ�`z��=��`N����r�3{��v�8�?����������e���"{���ä���}*�$���,_`����:�����Č�w?YÅ_���2qg�9� �x�a��u@�^��P��_�:�px�-�9�k!E�@��Ҳ� ���)@(��~S�n~k)+vz���7^�w�%��.=�����e}�����*~�˭Ĥ�����xL;I0_��?��2�����?Xi5�t3��oو;��%����P�&��]���T�	c�ȧ-"�R2����)@�/�fWu��W;�KI���A 3��G���ig�5�id���@e��R�D}x^GFfs$�] q����oX�ک�r�!;� �H��r
���L�SN�dO@���BT��i(�q�om�(ܿ�:)����+�IN�y ���J��+޾�YX����ߐ��LBY�n5��HS���0�*'��B�O;:G�6������X�ݑߑS%W�eG�R`�m����~G������<"�	��ۢH�¡Z��K���_��'�u��N�8�]�$t�V�G�Χu�ե�`K7��b���?�w���>����`納eV$�nۅo��
9�ǳ���3�Yb����� �G�U�YZ�Z��L:\�	�a���h�׹�.��Ad	�����F�ͭT�o��Mt��T���.�ӇT��kF����@����ӹ
n���IH��(�m��B��
ęv�F�~���s+��!��Q�]n��9#�p��e�Ν����bfؿ�dok����.!V��5��w��iȁ�}ЀV�d�{-�dx��ZQk���7���rɎ�~���ʦ���r�'<=����6�у�8���f��b�+��bB�q��b�}`����.�C���q݃�]Q��4(a��?�	���6�ѕ�W����,��a��_Lr/Ɉ�fj�'([�b�w�?�H*P|(����2'��[��`6H���}���lt�(�j'xk��������p0�m���_�sծ�j0zl~�f��5�O��!�_�"��W����~wdʯ-?D����*��7��+�ݫ_cGK�L|nJ����mZ(�~x�Z�q�_���dC��רՒ��BȀ<�-��8�����M�(0�Wvt( Y;s�x�ǯ�T��M.�\<K*yg�3Ft�\�]%jM �}�}�r����1�!4Z�]��~:��}���@�G�k#��'k�:�+��/
�F��s��+A�đ���)V�Ȍ-޳i��,3�Q7}u���R��K���fki�q�+�;���/Dù��ӭ
����k �r��ĸ�ۛC������z����(	��#ߪN� �J�j���,vP��y"�'��F8�o	�'����j�B�'��]͞���zjK��ۻ�?��?��R9?�`�
��1���[�e���q7J�<��S��5��8�f[�	�����n���i�	���!�C[�����=�w~����v�UWU㙳F�#o�Ӷ���9��Br����8۶�;k�� M�H�m�M����Y�H�����ύ�<�z��,q�ly[�
���Uw��1h^jJ[=B��.�3>t��+���ZD�Սs�$%���$�Z���as!������?9!8�������V���tE=�����葚�3mu&)�L�^;�	]�x�n�qDw��
��?���?�$�e��.��?�PO��#��v�{�P��xb�Ƌ�l���M���+�q���H��0x*xUQ*��/)��;�T�y��f�"���ӄ�o���ߍ)�u �[�
�K3��=�?���/�XY��O+4s��D��-�1p	�5���Q�	������}<e�'%���襐�%�6AHO&�Lढ़�3XjK�5��=[���WE���w���-��Z3����4�_>�̅�)w�{3��3�W��Խt[xq��w�o��F�Mܚ*BvS_"�Ś��{���S�YuI�� kP� ����,
?�/k1y�ߤֹ�(s���*+��
�9{B"�,o�/�Ǩ���g�Y\��N�?��P��D��u�d�*�u��:�8�eD����������M��5$����p?n�E��k�m:ϩ�dt!�@W��A���NeM�.�e-%��/q���P�ֆ\����˧��LL��M�<��r�	1�+�
��sYH%�𠝬�ě(��Qz�S[��y�O���v7$k�V�1)����+k~��3�����F%���^'�l��mG�Lm=�wS���w������?^���~���9��i����~�ӛy����g�>������I)Ol%��PE2�<�y�"{������
o��h�)Ϟ�f�eXwe�bOz�q�dD�7�����ձo)X� ��"��Z�I�)c�ű4%�]��L92����I6��S�'h�#��Wu{?d����x���}���"�V��b���|u��q�{�*��43)k�~����7�XӃ���Ǖ@_v�g����Ș$)���Թ ��y��S��y�����H��E��j����b4��dSB�T�)��ra���3&;eV�����]66���ڰ���7LR_Qu�r�d���H��>�k�(���	S��K�P����sM�eØ�Y��؈��0������x��l���.�G� ����"9&?�М��BQ(JF>�"���H�H��X�������c�Ŋ�c�Z�E�jx�fXfe=�z��J�a'��4=��������F���nq�ter?A��@��]Y�Pڄi>p(NQ���r5^�0�Y G����F�7��ER�ldwWx�I�Xf�jɼ�R��8J�����֗��� �@3�f�/S4�@%;��q=�)�b[��\0/}fl	�C���<��_/���[B�6w��B瓀�re�CлSN���
ū�0;M�H�9A81���J�xC��	l���,�Q��)Sb�Αjm�1:�Y16t���;�'�+{ҿ�δ���C�
H.~�u�r�T.���o^���v=�_(Is/8�2�/��bM�J���S
d{Ō���:(�����k����2�������:x�؜��f�q!2d����RpL�����?ʶ��'��ȟ�l���/�Ԋ�5����\C|d��!���'���7�J��s�$�u�T�hD"0&���Ⴕ\�4ӡ@��o|�t]�z��郪���D�}��C�~��;M���fMs㭉'���K���K̉u�Jy�qݰ�}a��T�]ΧZ����i]���s溔eɦ�3%jb0��PF�(�q
�'��E��c�U�{pt���#���J���Q3>:��]��-Zr�./r]Ug�G:���h��:cZ�.�H�w4����d�O�E�!�ҭ�O�۽y��3@ys�տ�݈]k���18l��Lh)�$I�$M��\����ӎ,L�MD�k�L�D��s�I�,1���^���I�eL���єm�q�n&0�i����D��|КW^#��;w����[��5>�L�uqn����Rk�q�ًVfM�rÃ�����!��mU��GZ�F�2�I51�Q�[�՞�G	�ݤ�6�.�,ݿ��|f��xA+��2�.yi�OT"�����9��S�����"ka����7�[4�au��(.2#7*�=D|�_��_��Ȧ��JnR�DS�u#��V��T�"�al�Q��Y����w����vҿ��	o�]9)�]�5ɾ������/jdۙzT��c�~��V�����?�XT٢d�Ʊ����F|����vO�;ő�L�2)`��ɺa<#�Ơ���b/9���]Z����d�n<�Xф#,-���`g�l�b��p��"h����G]�T�ˊrn��Ib� rN��$�R�ed-{/Eq-�)��n9>Œ��g�cv�Y�8+a܁x�m��0O�{R^-�c�6_��T���Q��8�VP��9׽�dW{Q��o"�R�)����XR>ݎ6���VF�i�ؠ�ޔ�ui�{A�Ƌ�����z8�a%�\�����6������>*ϡ� $�L�����'2���k"s�����'꥾a���~9�.;Db���z���C���cc�W�ұ��Wg�90A2�C�"��	s�bQ}
�JÉ�8�U֖`J�ˀǓ�~.���B�0����@���zo���cC,�����yx���b�]e�T�$�Ie�������������S��h�|�H�O �Tz�fE8{��!��u)SON
���]b�*��_��[�i��>�ȸ�	�iomj�����(�IJ&{ҫ����ef>~��A�>���y7^,�`���GYަ&=�g�l�����x��z+������F�UspX{J�,9�ڃ�\ˡ���ɫ E)z�NX�*�n#��׷h��}3��ij �S���\3�"��_�b��KSE����0~rpؼﲿ3j������O��k���P@%�7����i뙫{���Q>KN��;ƴ�ٰ�4R���K����++�m��n�|bty*�	�֦��I���̘!"WX�.�G���Z�|������`�.)��ݡ�E�L��������V6�Z6M�76%�2�Ð>q�,U+�&�ʛ��	�pt�Ạ��z"o�^}-�PZ��"�Р;�&��v��2�рU!U��Ș�|S�o�/<��_6��0���*y���^r;��J��`��" g�J�dAGu2M:�܄+�ru��ۈ٩�8�~�|�����u��A�\�����9��g�#xs���>�ї�y���ʛw cƒ��Qa�(|H�1���G��&����U�\�<�Q |	����&kb?g��5z$ء����v�{��d� ���g<�!�+Rd&��0ܿ^�+�x*:2���#�}���*�Iо�+������V����KO�5���\�[�"�<.�1�Q6�-��wv���=�w�~<=����`��q�vV^��q~|ښ����J�Fn%�8�U�;^�=��5S2�%iU��'��_�����I"ҁK*�#�|+�J�|�����m�!֔̨�H �n�h>�������j%���y4a��բ��v��A[U-���y�5��52�*+�S�3���tȋP`��,�yXƭ��'^�"J�@��UG�3�=�b-�TFp��x{��J8T�J��b�!�A%�V��QZ8,VYj�v� �t���Yo���0������s���m	��JB�uZ3{P6nM_Ւ�aG�*��
�.���wP`�ϵ��/rA�5���h�5�0~מT�hY��:�z����탩��0��Z֣u��$F�*#��?=0�oR�G��P�	v`����WB�5^؛�a.ݴ1���gSz��ҋWܒ��{U��|�1G�Մ�>�G�/��}F/_
��O2;,����૳e��q��=��(����&����i�NA����_/��A�0�2fª �^w,�������P���9��M�X�C�)M6�?@TCR�;!����H�$"_�)�E��]������a��(F�UgV��v�4����1�h�Б5�/���e�n�MT���4C&j����;�Y�����7�����J����AR�����B�G���*0ǂ����8}����̾���ಁ�� ��8Zg<�=�P#�R���y���w�~3��O_��.��M��4>�	{)�c�@זS�K\����W�X��8�x��2߼g�T����NtV~���ن�;�R�&ɤ�Q$�o�
�$�hy3D>a ��x}h]!
��GJ�b���n{�'y;���1�]t�+V����}��~Ҷ,���(�*�淿HB���D��sT�!׽.���YR]s@��t�b�;�)�����9[�7�0���{o /�q����}T��Xř�@r�����:ᛕ�� ���#��3���6��C��/�&�[�c���++v2F\�R8=�J��`�G��ҁ��e���Z�?03գ!A��-��]y^��6�ݜXPܱ']z�^)��"��M�cT���%��C��Fqb��,
���k&J����1�YL�݆)��,�8beH"��{4/[l�Ҙ����E���wmj�*����aaU�j�f�'`�ՅVAJ��q���%!�������4��P���C ���(���'M\BI�G$ؔ[��d�ځ%y
����!�ִe���ؐ��Q�Se���-Au
`�Ӿ)׎e1���k�(���v�N�V�k-��W�m��R/���������s�'O����z&���
'�p���V$��i`�//6<`�?�4F"PK�R�Qx�B�J�k�\�l�d�}:qe�A�; ^?n5}�g�H�iCi��� ��UsL�b:��&�*u�dJ���N�zp^i�"������B�|�"/\1<�!a6QG�K� ���u����|z���9�Ƭt+!�� ��U�ݪ'������x����������*�s��fe�5�ᦖ�y�ݼ�r*l+���V}d��f+'k\�;��gt�6q"�M���7.`4�p�"Ƴ�C׉��$CǨ@��$���q�Y0� ���쭷�pM��trzM��oE�^qi�U�/�Tn�Og.w3��T��/�c�q=b���Mg"����ϲ��i�d�2$��W�BEQ�ܱl=T�h�CT�箚�g)�+��F˴5)Y*�����[�fC��)�s�y��"x?^��k7��ԱS�����*�z�o�S��� �h��X��;5�Bn����TDG�����M�
�+�_�G];rtmV�~o�yh���0:�PT&3XU�їMG�۱W��!�Q�a�[Y�]bTSI��FU������#H�,�ޡӀkUet�H`,�9�zD�����43�_�J�K���rR,�g1H��֚��L��4�*��������참3GWU>��3�N��3�ז
\�m�`�s����g֝XAX	b�	�3�lm�c
����)���ov�T����\���֟�?��v�8J��b�s;�QT�l>�E����j��K]���s�t*s?p��Z�����6k�	�u���i@����>S�9�I�G��q���MU��ZLת=��,���p�6Y�ι梄���Em�P����/�*��=�{����oh4�M���`9�G���k�ạ����Ko~� ����]�"aS�ŵ0Y��QƟ���r��i_�ˍ��~i@QWK�����<9�@�
|���>7c��<�'@��A3�b�ʯԟ�l���k��r�aG����R͂C�mq�q�q��K�U�Pc��U6v��mo៤��`�?i@�j��|+���D�y�w�rtgE��8� {�ᣰ��G3O�T�Yq�=�+.1����4�����
c2!s���~�����}<�V�D{t��M�"�̳��ID>y�O5^�V�)��l$k+)5Z�p*�æwHcl(��ݟ���z��ȁ��ؤ
,�N8�F�S3y��\��SX ��%O����ǧ=�����&����K�l����V0T��_�r;VԬ"ȴ,y8��6��fiUQ��7\zvaC|����g�r+�u�Q_�����ώҨFa���℆������/�P��2�Foظ���9�?}]�u: ���aW��v��>�1�uF^�����)0�n�s)ĕM1 ���7o��hV0��܊���3|����\|���Ђ���c�Sb	�8�+2���z���m�P��扴�a�{�d��U㤈�%ʌ8°#�Q�^�����S���*��5`ᠧ�~N��ᠧ	k�7�!���D7N]n�\.�H�+�r�T�gz'6t{�ut����)>��%�����h��|R�5|;'luX慜��5��8��'�-�?VY�H��%�i�OTD�N�k��������.�.�Y�͹  ,0Zay�1+���{�y�{�/&$aYB5���
���d̹��#��2�I��°L���>Z9�Y�9vi��|�:Ww�mm�F���o�Q��8+��;d�ӧ�Eљ�� �n��[ �%ی���Pm��3Y`�AN��xn�>����������q3�j�2�aHI Y��9V��(���xiv0�6�g*K?�"��⮐����$�R(���RH�$B�����2�o�Q�(�i�$��`C�!�>�hFO"!*���(�M���E>O�:��������ߗ}f^(�]>�;Մ��)ɩ�VK��PK   ���XF1��^$ �B /   images/efd6e310-ffe8-4178-823b-653710540121.png\�\U[۽��n�R�S@i�n�;�KBP���n�M��tI��%�H��z��=�y?G��^k�9�{�k�5	SQ��D#E��`��2�j0��i���W|�~�\�e5P�_�P�gT']W��;���FC�%��+7uGK7O���'�����������Uھ)�&+�R��˟_�:�3ȇ��i(:��O�I_JvS���#���!�"�c��p��?�FXyB��%������V������_�/27SL<>�{n``j`���"� =l�,�B@ �a�7�=����3�h�D}�#���{��vsqO�����&��~�W����" �Q�|h�aV ��5Z;n �ޟi�=,م���ˠ������k��a��^�Ob��Pbq�d_Y`f���ۍ�}Q�3�t%�����Q��0ʛJ�P����,�+B����b�,� >�B�+َ���j���"b(',���ME$��/ف�ˈTt�3��`�x�%�J(�>]il�+F,gف�������]L<�P#fȿW�0a��!:=j_b�kH���T�G���N
�����r�^�����~�,�[��.���	��g����_��������ɘ���bǸ�4��n�f�;�����D<��a��qqS��m��t�3�0�YV� w9�����}�H4�:Ćg�<<0�������U���	����,!�1����9z�9�u�&�ؓ�~��9��k�t 1,΅Gɫ\/.+P�i�V�t��5��[�! V� ��P�jG�o�.lޕ忮F���"�v���5�U���\L�鿾(�C�N�v��t�V�Dĭv�'�u;�e�bà��<S0(T�J�����2t��8h��U�.lc����H^���~����KH�i	�AhY}N؁�0���0��mG���͎`��;2F#�����#��
0��x��enw��nL#����@�Dj��U�b'[$`I�,�JĖAU͙:lW,�XU6�"f;-L�l��,�W�����W�)$���89$��I���.�gJ�p�1�����l�N�%"�bgQ��5��Â���\1���	��s�Or���MMM���2�����aqs��0� �f��:���p�xʑ�?$&�����!���%��v�����i�FFE���c��~���RR�:>9Q����y&%��$ejJ����CE39��y����KK�����}�>S)TJ�h��"033;�򵶱y�����\<'%%C%J�Ɔy��&mk���2���غ��������5`TK��И3�9��?ف>S��j�g0��ѯ�###��=���~. б�H�������0�����jo��������oh6����ȡU�h��������l��`'7���j�T�7���d==i�n�hA2rrD�k��B^����]WZ��(��̾D�� ��mĒ$qss������x�������p�D���9�R�c�g�������m��W�Ķ}z�\^)_�D���>����O.����iˍڢ�=�EE3w+���a�X���x�	i�r��38u[;;9~ϷF����Z޺���R�~����o��$b��'/#��G2WR��|`7h�z�����cq1��S8��(���b���.%et�v5G�n��)^�X��C�c�J�ZYh����"�);ff�(=J5�_��t����	�����o�����v��˛�!�Nqr����x����]702��v���3"V��mA�*X��6�
X$���D��:���nk����޾����ǏM�>�/�>��"~+�}�'�����T�1J�/%$>�~b���XyB)�n��y� �1k 9�ct���0}djlbN���鏏0�;����������9�YK��O/��edPz�n�������'Yjj�~�Ʋ�b�h�22(9���X҆��[H�μ��V��v��m�3(G�z������mK�T�s�АB``��Ϻ7�K��X���h�+�H
AB$d���V��e�ת���p3d,J!�Լܼ�F�j����Aվ.ӫ�I�2�4n�m�h}�{@��#�n7�N.����*��b �!���$A���*�,V���q>����Bcu��5�#N�v-0o빁>���y���<�	������2]��J�����J�do���l�`f���H"�N&�w GDBR͕�79����;�J}y���ݭBS�+@��y�'נ�����
|:���6�,RM�{C
���<+���5�t��GA�}'
�d��1��Ќ����tvv�my�㱿��\t�� si�
��B���hׅ�h��c� ��(Z���V���GGG�䨩�-��C����������1bjzzTN5|�	
�����"\�P�BGO�߆�&7����հ����׊���6��� �|"���f��l�ش��t�q�> q��/�u !!�	�ddf��="%%5�C�b`�#�蘩�v�����j��&�d�AZ��z��ٯ&�˳#	ԥ4��eU �C<k!W@�$�SǱ����bu.�k7bRR<	gg�Q�hdl��@V�.����~�iiJ���zdlk~}��k3Q �`n.99��o(��tY�p.���>���8����,OO�X�##1�����D�:C����h�z{i^���w���j��yE���kRP,�����j���r��`��Z�����A���Y43�޻@W�¥e�~E�юMO���~>��m����|����a��}h(�B�3����
9���J8�}I	���},�3(ҍh���?�48=RQZu�/[&��ٓ4�m猟�,~�ixw+ ��yw����Ky9{*�]0ߛ�,�4>'wwͷ��LL�,��]@=Utt��]�������e^M"���r§��2����N���c��F���K�HE���ϻ�9�KM �u�_Э��A:�+�q��8_e�7;�|�d#W*���~S�����:�	YR<[��-,[�1<<�L.
D06:k��Q8e��x^#'��cRR��a���|Z<a�s����Ϋ��${l0d����*Rvc9A����t�ؔB8lF��k���x(���8$&&���z��%$^566��_(*+)�p��+/�:P�g���ͳ��2�TQ��-`�r�Ù��lh������5���=-�111c����63�	_IK��.i��uttHzxx��.Y3�Z� \�"�K;�w=�ē�"4<""������Jw�1z�\�����>=͙(T�8>>��s\��I�[����k�װ��Մ�[i��-UեV�W���_���@����fP����v�M��������NP�z���'�a1���Z�R�p
k�
���M�������x���Uyf;�8L9�-(��E8@���~��=�(�گ�
���zc��w.����aS��OL��\����Z�aӫ���?��QPx�~��~��)>%T��a�lErBS,G��Ы�9�!�K���x�'���o؇�_̭��"���d�`**��.�*N�ў<Wa}�2Q(�{��A�ЋSL}��p��<G�=V\\��j����H�1��5�%6��z�������%
*�w�#��GfӽI@�IO�j�JJ�db���k;�u��\]ёEn��^w���}�0:>�����'�"�B ��L�уG�V�ϕƔ\���ܟL�-4.�����iC|߻����D����3��K\��?��p��zwf�w�:k�q#�NML�a�4H�d۝�b��M�ScZ*ʮ]�2a��5��I��������Y��u!�/������ׯ��;=)P��BF>���4ܵ5��^�p8��WEE_?2�È�YAJ
������y ��@I���Ã�9)c���K��t��lo��^���F����Z���+����L��cQ�y1�h�2�㇉��


������v|�b�Qg2L_�J��\D�:=;;��XB�UUU9�=��R�PZV6V�F�ٛ���}��bz%LL����MN-T�\���F����/:!C��O���۾����޵�oj����3����h�,��쬘�:> ž��.��8��}.����x��	[��,j�f���ހ0�]�Ȉ
|���6>(���3��&wt~�EI[ۯ�+���!!����-,���^�pd�>���L�\�G�����j+��zǑ�Y����M�N+]��		�D���w'%��������ݓNM~l��;u��*/�����ݒ_���(�󕃖��SjFP}?�e|�B^˷o�J��0�����������?,¬��x�V�J�`�� uT��-f���,����/�R�W�ëPz#1�3�R�?9-��c��ѵ@i��렠n����G���7�xxKO���Y�4�=�3wxtdr�����������Z��W�n����,�_M�Q�7O����@J������e��PIj�����:���<<e2@��miiq:Zy%u�������21:�c������h�.�O�ψ�p\����i�?'~��\��>KP\N�.uw?�*������L(��ss$��C���<�H��9�}L�\}bphT��~����CR>����X���k����"Ɔ��"��1==2��.���P�c| �`�? Y�	����r��.���B�ff��w~�N`��w�~ ��gP
lkk�Q�{LD�:�/���Փ-�U+��`��0I���l&�( L�S麩f��:Vf���g�8�G���N�n������~6M0S�?۲-�шQ�����P�w��X�]� }��^��<'?OpP
���d��ʝ��.��oWZ޳%���<��n6���ɯ��Ѓ�3��8��@ �Z��w+C�vFP=L��A�vw�Y�X��A��f�\���Ҩ@u�I`��ku#�(O'֎U���Φ��2����襄�G�^���|>bG�;~�<�8���/V!��J�.@�5�!���Ǌ� #7{��W����K������yx��~��� 0��-�@��7�s%M����]��_����Fm��s�`��y,1J6y89ہ>p��r�<L�j�:BħW��!.9��v�E ������'�H�4����Β����g;A��e��{cD�BA,���x��.��O������ⷴ�.��p�Z�fܘ��a}]��s�l�$B|ӵ��JRRn�J>+뉐���>h�#���������vV�m���eh�i>�6������o>Y<�\"�Q�֖�t��Ĕ�g)Bkc��뺂"+ꩇ��~}7��D��D��cp�Cz&V}	$`e�ӭ�dA����q@}����N��"8} (ǧA�,��95���3�(�	H(hh�l�7~�����=,���K�z0ٌg(�P��v�%16�=?���#�.
9f�(sh�����U������< ��ُ����cc�Q/Hx,��v���୉��(������e��>�խE$  �*V/�yA�9���Bc�R�'(���0�t \�]a�x��΃\xYkx
8�AO%�b�<�8 �X�QR�9t!�*1Y(g9�L�~cN���'`�t\��t^y �ֽ�ȂvA(Շ�6Q�uA���%���)Y���lbAք��8 ��K#�YY0 �RNN�C���d����vKi�"~׿@�FJ7L _|���90�p$I��,�;�h��3ZL/M6��Q`��(I��U<F=?6�ڤ��Ǥ�k��=��W�U�TN�� �	^�i4F��0�U�f|��������6o��SZ���{]��ˣU뱜�,����fW��uoȎ����|b𱫱��ay$j���b��]������ojJk�����A�֖`��͠�/�uP!w�uIb������-	���`��E 1���% )���N*��6:P�,��	N,����n�]LN��7���l��h����p���s���g绛� �I0>�@K�L��� � m���}y���W�����v� ��J�	���
CaI)�C፜��<ڛ�Q��c:@�Ʀ�����5�c�+V����*E��Ӿ�6���Bs�3Œ�kjg2Y{G�xi&�����0^�i����J�L�n���))aCC
���Y��+�륁���0���<*B7E�gA�����ɠ٣�%x�4~ǻ� pi��wо 0`p1Taa��m�׵��O��QQQ�&��N�C z)e�JHH��[YZ���4�{�stf&$(�a������/O��G��x,� 	̏�J����D;
�(�h@������������ё��4K6�I@�*��龣Q�[\;Ss�9b������*�z�%4Y_��t@ڞ�+���6A�8�!--�Β��]��KG@���s�V<�E�3�D���a���Lt��`�e�O,��m�ڇD����aQ���Ƶ���VZ�P��T�e�����Xϵ<muC��M�8R���_sj/yKѧ�|ħ�imm�mp�]�y$�n�L��*IF�"����#�����K��������aa&��O%��o��"9�ఞ�J��_��&�dft�c��V�*��)A$$BKI�cK�����@z�2�~�� C�I���Ǿ3UB-AxH_���㰰0#CA4tt��a$����_��� =0��Gqtʗr t�(P쌥��m]|����jOT�j��S!!!�b'}I�|��tP���æ넉lz����y��C[� T#2.߉.]�����O��5����w�q.1�9
4�׵�\����]�'��2�;�_���<{�����all300 &!�><����a�� �2�4Zn ب����C��D6�ϵccc:��/�2E,o�YXX ���|��/o���9�63���0EEŞ7���:�l���q@h��O��f^�.Sa�V��5䍙�GP��"�-����v� ��� J"!cu}x�N;}o���D��ZÁ<������{���=���	Ļ�xM�����ѕ�k�� ��� /�[��\SwQ ��D^^�n��PmԎ��y�LvXh�>�a�y$�H5�ޡci��]5`	=��1�aK��D��rg�K��f�|�B����l'��A���k��&��7�WOfFG�TTp��u�����*S��^�-�C��dBBBr%B�L�����O�'������0�D�h	j�)))�V[ � yz#�J�����F�%x�����:��R�"~l�����f =??w˖�J����z{p��.���g@x��G&�=�E��r��P(g�{�Z�)����SS		jo�|=	����t^�~7W������1���n�Ԕm����E�����	{���6�^q��)gq/�w`��76�3�@U���u܂��L@�]j���<1sy�`���� ������)H�P��4�3�k5{��2�7�3Ӆ��mu��ۋ���D�h۰�q�2�J����j�;%]����'S*�Ã�޺D��	���`�>��v>���	�Upۙ�-���!Cʔz�LG���(�A�K@nnn����!B�VYh���ق���Zl�9��AA�{���xp�'3���a�'��h'�tdf�u��{ &�~,'��p����/4�.�upμ�p�w�.o�Et�[�����Y���Cū��B��te®�{[�$����kN�^��Ƈ�-g�*�_7�R���������in��K� ?e���t`sz:E��R����u:��*�^����]�^�]��=�qy����V"�(\� �����wI}uw�Ly�uK>�tl�hr�ݟ-o�u�Y��� f�A�pD��� ;3����jd�2?��H��k�_����e�Z9^�3""bye��,R������Xk;�אV{uK�u���������A���I�ίTmmmu*����rb�u|LI!�������0j��Y=������v���cYY��=��J���1<�X�����V�殔�*�c}P^ �C�|m�m��y��0$����߉܊V�xAPJ�0
��ok�,��z���,��)�̣f��;n+F2R���L3�/}�	�0o� -�\����Ǐu�X���|Szi�n������WOƲbQ��00�����k��C��"�ﾫ�����߆�'X���y��(��Tk7Su|*��^9c�]�Xf %b��:���q����)ٞ���w"�:*a��XXX.t?kk��f��$r`��>�`�c�{����������Ď�o��ã���w��$����I�##��Ρ.�ޭ���1�?�Z]�р%<��\YATWO}�:gmm���b5��p,mP����r�С���	,�F�kA��2�N �|;_cC�h�,G�������s����V@]]��nF�� �w�?#+k|��̌vyr���c藌�hh�ڀRR"lfcd�r�ܝƼ8X��yA��D,��мa�G�~�G�9H$��/��^�mn�M�����,��<s\����W������m���J�JB���S	�.]MJ��X�������Bt���((��B��͂��C`����Ĕ�� �tmY�����t/�\��1�}����A�L��`�^��!�?q�#�+�>I�/-ο~��/���Z���'xa�>�ss��G.6/_�|�O<�1�<�,�r�;�k4��@6�oZ�p�KL�g�@qI���	��b@4�*#/�y[�����ܽ;5��3�S����z[ҽs����$�k�Y�)����y��X��X��������P��7�2���#W��%%%������(c�~H�����W�2(wvt�#!!�Ĉ=1:��ڤ�:.cŦ1��`L�����g�ps�i�߮����oSk3{���ѩ��m�l�ӡ�"����l����ފ�C둖�D�2b�������b���GR�8_���n�v)���z3|����'R�#ss)	��UxhA����VVV���|E@��?~��.��8`�¨o5�N���}�9���{�� ��݃2xFRW��炚�Y�4fd���%!)��4�(���M��f��UTq��u��#mZ<�����PA`:9:Wd�zm4�:���j����z|��o��zG���ܫ����~ G�ޠ9&<�e�n$���2(�,��&	��\/R%Q �6BCc�rO��le��꟥6�%��_Is����'<{7t��`-�u�o-�?K&�bD]|���;ƾ�:����i�����ֱv��k�$|P�am���^�kN<��6��R;�$���	H��CGG�/�`k�]{\���B�����| X&dh���m��Y�$�T��^��}1�)\�a������g��Yot®��Z�F����Օ��ޮ�������h������� �D��+-� ������� �-����]�)��q��������'8(]�*�1T�r_0�����Z޽J9S�sWi7�c4�w7^RWZe�!P�=���j�('+��S]�3�
V�������1��E������V�(1?Yz![\ClUDT���
_��n���Φ��te$�NJ�O�KrP����Deb9�hq3,*����P�rQĬ\m���dCQ���
-� ��W3�+5��-����EYY
����#�#CC]���N��_�D����F�%�(&�X-dc��m=^Dy�w�ث�j���)�!����݋�|����<1 ���ab�nL���/�7FHHX�W������7�jۢ�u���:�us��/;;�T���oc�_���bRFoAP���a����ϱב������.USӑ �i��p�=�(C�q�vϮ��=?O
��L�;���r�o� �u.,�p��sx�v;2���+������໻ޭ�]j���I����Ț�������Kgh��u-5��U� ���P�<s��AQSS���^S�,/?�G�O�9��ַ{缤��]���i
�����*�]_5Ktb�N6�we�/?~���]��xx1�\�u� +jmllBCC�$% �=�1R���'��U�A�ZT�
��Q� H^hQ�����a�!عV#hQ�����4R}7"&���¿L�2�7,&��>Tx�Ը��o���8��M�..���d��n�f�VYD,\��Y�uk��,��l�ѓ�q}Q�9�%�'��TI|���O�T�m2��z�1c�������#�/�1y=St#��E@��L��T)�-hA��T�AZ���Y�<Z%~f��R-��4��j����|�����I�;��h0]<�n��d">�
��nZZ�C?~�J't]�O%�6�"��(z���͍���`�NI^�cJJ����G�8��4|��檿L)�sq�����x��JgQ]Y)&.�AG6���9���P*o��F(.M��H����)(�da>�khk�m�x�j�Y�d��7⿜ Q ��R˼�]|V[ä^`��i�W��~m9^
�,2N����x�D|������=i8���;N���=������|����+�������Z�5n��P?{�<g�O��B����He����3ԑ:%�`$Gun��5^�w��� �@�#��#���Q PW�Һ�dg	��a�~�eE�|lf����@;�������1��+)*��ج�2��������G��uD��nA/5�Fjhh��kw�q�����BN�Z(0�:� '*!��v�6��{�\M�����.��]\]׿�)�O�����a�n�θ�||�G�� vZ��Bp`�Rȫ]�u��p���삎nh�g�-�ۋ��y�A��DDDa$�����}�����NN���&ê��/��v�����Wp����=@�hx{B����uR�`$������OQ��'R��q|sX0\\\ee��j8�;�I3�N� �<���Ru;U�m=S����!��1���}a�6!��EW��(����}A��F�q��v�xvv�m1�0ʠ��ȝ�Ҳf
�x �6��q_��ݧ�WwV �wd�����\�v�q���p�\��7������[�ƳYX�/��w���ΜA0� �@�U�Tl�'�ȩ8p��kjjj���)N�@-���Zu��n��M�`caY���5����C�����>���\��q��KmF+~��z"Ir#+�6O��@R���Ef��`����ا���8�����tRH`� 	R�x�!����=}�-�%F����j�~�٩�YܑL�^ x��bj�֠���_���d����8-1����~�6�F�����Ԯ..���1�N�L>|8[c��ۦ���u}�R�X�r}slx��Tll�4�7k��mw�)nS�p����)�k��۲�X-���ק�����ft�78�	R�IǃF�ݭ�'�AJ���E8�|���Pθ<��E��?P�<��,��X����ݶ>M�N��o!��9����Ea���Zg	C��j��Rq��{w�b<y�Q_�T�����q"^Z.;;;:m�s��P��q%(��K5&�,���Lf��?������.>~�N����+V�:��M���TR�a]ה`�?b(�Õ3E�΢Hy�HI����A[�|F�\7�2D���?��p��c!Ϊ��{P��Ok�����4�>x~~����1�Qk$p>0F����'x?rTP��U/��1��@�2o�Y������w��o�P���'�/�Y��y=����Ƈ�C'���@���;S�����DF��1R���-��/f�@y@�O�9���e��[�ب���?D���.�;2!a��=�����4�ќ��j�c�GN��_���ë�*#�뛁H�����W�C~~~!�K������Y$=��
���8,�!a`�ٺX��cK5Y��q�T
F�d��z��t��U``�F�����|��(J���l�^��E�E��.��lkF�wfV)Zv��D�@��WnnϠ��I���G/@�WTTL���������ǻ;�	
��n:�jښ*IR[��5<�Ţ]n~:��+o��!�ϱ�(s��D6���G�RQ�ra1�l,,�ت�� {@�ko~�-
���f�r����I�ϧ˭ 7�����r=�,K$Һ(�����<Ռ���pyu�#`����&�����1����y��+95.;�U���>_h-*Be�m�d�ae�5Yf�������2w�d^���3���E����g�����h�����{�����y�X�(��jJ��G�A/��`��1���?��P�,: TE�\�@��t�ǰU������$����޽��p����#l����g�����N�Iz���E+����ڙd277=;;X����)�^��
��{o/2hS_��m�n9�~�%8�i��$$ HH�|��꼡�Hn�F$%	y�!�RG�5���6��O�\����#���L�NfF%h��xb�+S3��*y���_����7�
ŝm���N�[���C"�}cmc�����v��AjJJq|r���2)������W������~öwQ�<V��?��Z�C@@�����u�3�b������2�O��ٳgЁ�F�����ó��&C�d7�����w�	��b"��~�lIw�ar��o~�
I�������׵�t3Gh�p0��K�4���j4�d-,8�����w��2Va$Z�O�_��{V��')������ѩCD�꯬�_f`��Q?N��A�Q��'�<�b}�5$F9 ��Gq�<&��ަ���۟����H���,>{b;����vX��A���O�a)�?_���<����	���:��z��/###rþ8�p��H2��͕��N�62��~�炡�|z�������tt�~5����OOO'�冎�q����R�;f18G��s�D-�_�,+������t�@%o�)## g�^��{K&6Y��p@^ ��N����������;C@{��A{�%%,yMm&�
dK�H��A���\,�=�l�Nu������뫽1�''���� ���a###7FkB@������|C�0�u&�����5�F�BP�O�].#��rN.�K {�T�(�����Ѫ��]ׯ���ez�R��-��d<���:Of��� 3����:G�bO�����\��I<|�|Y�hP�ѵkɵ������wH�z�`����9�:$C�}i)3��?�b��NO�O��+(��G*��Œ����,*�w�����h�<ZC/ � W���*��VS]�n-!�UGg'����N�%&�Iډ#�v�[`��NX��d�G��$<sfba�g��STk��i���kKj!�b�	�9V����v:��v��z�7We+�/?{2���g��! @����us	׸p �n�%�Y*�߉>!�<�0b�'���8�Jl &����ݶ�����+++���Y4�ar�!ؿ����UI��̾��S�ܔx�+m˥�pOvb���5�z#�Y��O��A��3*&&���*�}�
\�'�7ϔ���A4����)'55"�C����tb����s0^�ka:F�RQ� ��L� � `Vm{���А��+����Si�I\�u}}�����#LҮ�F�	����))+���X�	x,��E��}���T{)�(k���/_�O��$v��C}��ɉ��{�)>��Iā�����NX�>X�d^;Br

����Oii%w����@�T���ˮ�����X��"Y��%�I=34������S��ÓE�ERy����`P<FƦ���,���m�T[���S^�@���7F���B�3Sa$��]_�,�̀��|���'5ݶ��*�8_/���!Z�P�. E�N��Yu�o�Is���>P"2f��Cv�ۜ��m��SYɊ�j���б=�8���jojJ-$$�&g{�%�g�Ĭ�@����U���n�<�Y�����_���`ZR�����}�-� ��SJ��5�x}O��ަ�l��KQ=H�4�N����X�Y󟯱A��J�`�*���}���OBJj��PڍSRR���&X����L�;�3�@��/9�P�@=�F��u���?sH����ezDXXX�ES�̮����PQ+�,��s�a'���k��=�c�W&��e�q����<TR���:Q"���e0�b�NN�J��ϰbz;j�!�]Q���Z�f�99����Nu���FR���ۀ;�:��w˴�ޏ��3�poT����}`kk�MU�U�~�E�n�+b)���RRI�����g;Tgg.��N[�O��οQ n)f�������5��x����g��Ņ:�=N�\@`�-c$m������^*��<pU����x���I�����r�>���\�i�$�,�`>{ZLY��I544�)>>�)r).--��G���Q�&����܏��R�,���W-�t�{?��@�
 �q����#��w<W�� `�x{mY�#��F�͞�Ϫ�8
��XV��@���lߙ*эH����[� W��"//o���I1����߂��]	,�y�%���NI5FA�x�����"�mZn�����-1� ssrs��m/��@��pxq���6�k��	h..��˚����h�����Iw ���� �ss��4���{��9�R���Kߝ��i��Չ1>6�;i��t�t�Q��g�~��>�K�v�̆�\�s�GY��c��p�u���0I蔁�����[��fO�Ko�*t��Ѵz�ٛ��yV�mB-{��W�f�y�c��r����lll4�UWSS�w0h의��˕^���Ѱmgq���9^��t��F���z���{�@����ɉj�E���6�����O�g^��`b��E��������VY%%���_�����~ק��f���� tFA��L


3����Y�[��$P�wmtR4�I�����I��~��J�$>&&Ԃ��r�dYc�32��V�i����߾z�N�)��آ�L��k(�n����;m�1�B�*����R�շ�}��`=u
��B���K���/zp�ᾟ]�d{�sk�z�ۣj\��7_^��}���!����8?�R�0Y���H���496CUۘ?ݶ�\�X�3ϱ�r1g���,arU7J�0�?���t"̎f
 �Jߴ˘kW
뷽30��\ ��^�L��v]$	�n����ק6pEEņ��5�z	�m���t?��p���@�� -jA������\]ɧ<n{xm�+��	|"� u,-Q���/���4ZFW�C��������
{����e2�gэspp���/+���gObV�߳ �0�=��DB"�O��(�/\h	9���Z	Z�,pP{����c��� �����W�v/��2�byT���8�ļ����@����1Y�U�U���j��7)L��8011�D�T��A"��]�/�-h������7>�b�-Ӎ<��Zv��Sh�@Ncb�x|ˡO�9O���%����	�����d�3'꟭�tCA3��`��o>��Q�����k����x0�p%\��-8~�#��T8���ƿD~
S�+�[P��/�J��	�?�dN������ٓ�f�����]ۻ�@�I�<��66���#�6���{�g���ڍ�]ü�������_!�,2�m9���� ���>�Ձ�>pߡu�> ck��:;"���SB�P�G3���.%��|�P�U�K�ho�
{\�ھM{|;���=\���!m�Hۍ�n��sEa~>��^�U������L�mE�'~�����,��n��S���~> 8��'���ߪ�q��Wb�7�
i�Cʚ��mNK�Ȉ�B��i���xm'?mA�M>"cӾ�: ԇ�B,k7�֌G��\g��xDӫ��K�3��������F�Y�"�~�X z��w�����'�( �MNK����#��c���I��R]|�Ka!�jݧO8�9��T4a ��A�g�	�-�����y�
Ä۔�}`� \�{w}�a��,����QN�iV�; $Ö��31c���g���#����{�ϝ�l����|i��˽8�������9B9Sdغ��s|ww��FW��p�W�{����݃@B����&�b��� �p쪦�ww���e
�F�{$�J�n���Tv���"�Qqq��|m���!��4N��E%��!�e��}((x��,8'g�� X�>��*5��|/9�ܶ?��T�|ϱddb�V�d(�ø̞�� mh7S�
X���>��d+�Ƌ����5��)K���U�6
oZ>|Y��!��UwJwww����!����ɭ�o���H���ٖE������fYe��4E;S*�x'��#���EBz��[@	B�/��h��#��}�����%ζ��p���n���|Ob��׃�>o~�Y�SR�O<J���W�[ϝIT0{I�ģ��		�oޘ��Ag��2E�ʱ�,w6�����L 3K��h�� �^s�k�Νɖr �K�wL���
恕�U�(D}x�n}.�
�I���#��[��;������d.���������P�2�����u�yM[q|KZ������ l@pYڀ��?<�G�XT�Z�z� }?�nm���@p��q	>��gggc�V�Rmy�*LLL��� .���0�^_Ԇ�����ۯ1ۤH�Q�=�Ѣ:��d��T�%^ا�t��[.�
�¬,���JFuFqUUggz��j�K_a�̊�r�щQ���������b3뢒��r��j�ꏘ��;υ7Ut.�$�cQ�z"�76����8�B�m+��u���x=<�%"���$&���T� ��Ca����C��IW�8ۗ���{'(�m�m�/}�������p�r�N����C{�ԡ.2Jn��&�����ko���k��(�g%jԆ���W�'�<^���ȃ�D��7{��m��0��^]�{L����5�T�-@���o������恊qr��9&u��;��7�R�'�#�@�o=��#�#2��
����"[���Sz��LNN���<��R�+��lhB��7|�D//��	,�v�����RUߊ�P>�+v�4K���?&�3��f����?�����>Md��adz9�롏�_ѓ+_��E
�-|e�x��uH���L�+�"#�n�+��¡o�<6w3q��F���rt[���}7�#z����ct`}��g;S���� ]��lB�J�4�����{�o��l�.�Ɛ@r��K��n <��߃6�_
����N:(�x����3.�"�u	f�l���?������2��g}%# ?�!*jp�R��u�y�WS7���1i~ڠĽF+Bo!�C#3������ʽ
T�Od}~m���"o�U��]�7�ZZ
���V֕35��t��	s2��t=���6��n�ӑJ��4иy�"]�����0�~�]�6��IȒh�Ɂk����]BCC�j�z�������h��*�����躢n�a��F��N��m۶�ƶ۶m۶ըM�}���1�{�$#�dc�9�5�<r��)}��9�Ƀ�`�������`��=��-==�ORJ�$ƨA��`I��M�iP&9�;�����kC{񇫔�F�X�V뤾�"��D���R����Wgx�� ��OV�,v�es�Y\����jM�[����xȜ�/K!%%%n���Դt��&~ C�
�>��jA�ōX_�~���.�ίX�/���mmcBBB����#'���54򊊊���Y�\a7}��J@���
����@�a���^��(XY��w�̸�踅b����b�7��
 U �s\���y/ m�ט�8�o�u}_�\G ���}�{8?;˫��r��G���s�����z"[~NY�H���!T�@ o�P�f\OoLMɛ~*��6m�����OV�Y!���<�m�)(�/!2����ꄊV	��%�;4ώ���g:�� Qpusk-vD�Gɮ#�J�@�S��irj*>-"�u���������00"�*��116����E�潇r�Fg����:���ݾ���L�
�# ɢo�߫'���ѐ���*4�#G~��,/�b��]]ş[%����NV�F��cY�g�9���A�|�����ni��>(;(���u�:h�f@ ����8����Q����_\x��B���� �)yG�� F�`֧��x�@�Y�3���7J�ǧ{́���F��?_W��OI�
���q�����_fF{Fk݆:=H�ڤ�q�������٬]o��,,Q��s�H(�~�"&������"���ZΠ��~��q�t]\\�w��ԧ�H,LL�	�GЮ1 ���3V���>�㿰h�gI����?��h���L���4!1qJ�.}��ǸD
9Wʒ3ď?3�3�6�U��-�<yX<<��� ���34tt��)�����������We]
`K+.<�����3�#�����E
jVDM}>�]߁��ohep�VK��{B�
�s�${vv���雙�\�{{����ʪD6k�"�\Ã��u�sn�H{'�fI�~@��$�i5�"��\��6�Vi a`Z�A<���![�ݪM���x/`7���` �GFN�܁�������	%2�����Z���O�
������u��2��~�q��6��k5_��S��HZo��g�z��GV�F����{����yQq�?j�>�����n��U�¾?���Z��B��Mf�����CH����_5�"6C�H��5�`��{v���j�PD�����J�#�qP7{��$�˖o��������2�����c]@X�=2X�'.YG{q)��:�h�o=YIߐ���\�v�?���������p���$b�7`�m��ܸ����x'���r'q�ȭܦ�p(q��n��ƺ�3d�d�ȡ~@�o�y��y��IKK3Z���XZY�Z�O� �XϏ�X�p��M�0t!N����6
�Yi���aj#�$�{,p�XA����	�'�����5a�a������+Ht��s���,8B�Y�U�x�Z�+������kV��9�!�<q������� C�~��KN��~-�C�c�����~� ��C����x=Q����	j����z�[�Z`��m]�b&���-��ޝ����#]=>�?i�C���L���4�WU66�~�ih>�g�crO��gI�+�*�)�e��pf4�۷�����b+Ɨ�h.qR��E�J�}� �u��\'���1/;��4P���.��`ڣ��xy,�&NP3J��������:u.��Z- H*Q �~�g7(Jhfcbn�l��j&�q�順^92���X�����������E}��X����b�~ x_d4��<�N6��0@��S���8��׫���rp`>#��Z��o��ํ[en.Xss3܅�(�Ƿk����1�
ж}KjV�փ@v9�l󦻪�b�8Qp�������FYL��㢪���e����C��Z�	\�]Ͽ�H7��F�Q�wv�v㵴� ���(�A�)Wbrrh�PD7Z@�a1�*�����8;;��E�ԋ����6��\]N�����|���D<"���ſ6-sj����' ��ZC��m)�lmn��"���T cc���o$���[����l�9�,@O#��j�u-��E���s�V�������C�]��d��G	������[{�SG_���0IX�w�� u�Țv9� �kb3nn~��e.�
���8��]Pݎ|�!C�����ˆ.� ��������5�&��|GYE�ofi&{��ݔx����L0w$�Sv�����$E����a���B�}��qqTr�}fS�v~{y��E���w�vS��Q���WGA[		���>x�?�QW���K=AG)e�4+r�Wjj8AAA��x��|#�}²F���Ǩ������~�ߜs۠=��k*x���;��K7/���Ƙ{�%Ʈk������m��� /[X�t�ܣG�;m�nnϮ#K��"��8�H"�C������|Zֺ��y�bw�r�0Ҵ�֬��'Mc���0rqq͊��U�,V����j�����pៀ͢���x{���Y��]8�l�FpH�>0��>�e|��L�����/�{�f/ɩ�F�ѼBYNNB���F� �ml���G�{;%�"�*FEMm`~�^LEݹW�P@0�z���V�[�\����WT�Y^N}zv�7;�\]]ڊL.�k���*O>,�Tl�z����;��6��M ��@Ϝ����'���	�֚�����I�Ȁ�|��\�֫oo�A�VH�"t  '�����tm��F!�����\�O�sb`.���	�%�P���qB��D���CE������!1t�$�]�G�D�vPF ��\\큍���ff�M�


��NR�44}'��%~7x00��=vVV����&z�<К2��H��׾B�Dd�_䩁n+���&#�-�
&>��C|�6;[����:�df0��Ξv�{��g�Pd�����5@L��$���в���?dRa��Ryj�I�h����]��R ��j�������C�%&�:�ʌ�X�N��)��������'���b^(��B$�h�`y]�����R�Bdp��h�.uv	��%z������Y�8���"?Ñ��րA��3� ����9�;	`�Or����ml�h��YO�^â�.YhII!N���<=� K���E�k;��Q ;�Q>��ǀV;����b�{���F�Ouɸ�p?>>�b���>v�>aF_^Z�J\FMNN�6�X�ͭ�ge���[[[#�~�&�2�e�O�Կ�Ծ�#G�κ��AP_0���}�v�ͻ_��:�}��z6����VIx='~�!�_ZU�9*��H����������sЖ!������r�>����III�qq]�8����@�5�wf�I�_|>�BDA�_1#�_�eM���CCB����Au:m�� 	��?w�&��f����#�P�p|�����y}m
T~�y�~v��ڮs�����c�E̶������	=��y���8j��R*'�>�ư'^9QpQH1ժ��y`��v$Ө��X�ϮUD��ң�����x�%��=�~I\��������Z�嶯��@W�����Gp���g�T`����x�8^)�B�\�:nB��b��;`�0�a�SY�)N���+��D��aA�g�Wb"ڶ���@��v�1��E��V55a �]x��B�D*C�mwAc����pGZNOO�j��0��%ύ��?��j[����I��C6�/Z�@ԅ*�IDD���NT���1�����80���.$TnQ��9b(����3�5%e/ gwǙv�}��
���GFJ��H}|@�SS���́W����t,��s��P:�����im����,�������!�&v��{�PD}P,G�L��
*c��MI��O��9�5�?�����m���T
	N�����eeLmD<�tXB9W�U@�o�f����n�,I��>�M�U� �b��gM�99�����<!��3�1h�P�c����T�6S�LD�����z�(쪳�"�i�2�ReM�����	A��o�}���R`���*ҿ ��&��\�mEZ�ݼrSC�]1?ςHM㮺���O�>���fBI��8g���(Q_w�������d ]J=�������(�K����������~s}aE�a���㓬{���vZ�_�5����n������K�8`ni�_�T���鹿X���E�yPQ�Zn�}��b������y����m����8�K^W7fwW2�� K��)�}�b1�VWWo��5�έ�bK ))�~)N��𽳳���#�g�$nƵ�MP�^n��kl}�_�o�$lt��.�s���:�>
�Ʈt�~����\7|�\��c*]���#8߭��3�ףݷ�l�H�ҏ}o���i��qE��oc^ސu�w����ϖ���������		Rnn<hx��I�H]���H�F�����{�w�zHz�]N�!�Zl�ʩN�Sk���l�ev�X;�B&.]�9>�q���
�o7Ya�Vk��=��������>��(/g��});B��(|�����DJ^�EX^UUt��[���G�H$� z&�t۟�f��IKnnn@�#�6(��iQ4:*ڨp�I����@��B�����jЉ|QDc����� ��>`�$��i��:�Ч�جW�sss]Gby#@�~�`�{4�i���_Z��$���1*�O�3�� �$�'??����q���Š�SsЦ:��3�ޏ��HG�����߿�VT�� $$&�z�A������-Wj��>y���P�|ff��vS�ݝ�^���!��)M�����X:
����^�L@U3??d/��<U�v0��� Lu�DAF�aOO�������ԥE�����t&�L���17Z�R9�7'��g��SI��U���2��D���f�p��*|O��oY_���	�1lZDL���=�vrr"##CN�-.& n��kVF�������9a>������T&f��A�ąr�D��bH	U���>�6I�l"�VT΍�]�ʨxl�9V��)ց�F�Iʰ#������eAU�I�b����yy
(�66{��`hhh@��vv��,.)�h.���}��Ϯ.�ɩ)@f����v|\����+7w���G[w`  -H�a{���b��l�ooϰ�z��G����)��������Hn>5������Z_�'o�;����+�6����ϟ�Ս��$ �١>b���o[�����C�AEg���k�G�D�Ԩ��<U�7�l[�:�X�$&��ۅm'�{V��V xG����8��{J��ŕ��k�B\_Ձ�A	�i�5�����M����PӍ��o�:���$w�J"����&'���cV��Zl�h��&D��/��Ӯ|?�e�Zi���ڇvZ
��	�����ۛ��3LJ���Q6WP��~&� L<��Ea/lȐGb���Z����X�+����}bm�>. δce��^b����N�����/As�Rm'��Hi��[ �
�C,�w0k�є}y�Ê��wo0���h �A���� �<,z�N�86xQ#R��,F'���y*���z͛*�����Z��񬄄�w�|~�֪�,i3�ŭILW����8����;:
+O�S
�G�ᡱH����B���7�=2��D��['��	��xm ��v�ڋuӒ2Z�O��DEMҎv~�&t����<=HGAa*�?�j����;��O:�OjP�C�Y�B�K�����v?�݂��:��4Y��묃�"7;��ӨH�՚?��56�~�,����0�ZTW'�h��米.���m�xN�P��^}��c�h��T	�8\�`��&;�Q���.כ�Lˈ�{��=��			�� ���l?~STS�bW�����4�Xe�����C�������u�;�Ml[[^s�N��y�Ux��t8���<����uu(}}}A'�YX@�}�T���3A�+^�xJQZX������uǽ�N�o��+��iP��Y�\I~}5�7���X=��ݽb5'��TcQY*�!��_&���B[�=��=t���>�d����YQ���X���)<�ι��~΂���k�4"�)�TߟY�Zr�}�N�;��gjPn�x}����u�<�Bd�B%�,1��>&nv]�٬C������n���"��8��4���xU�HKS����%]2WȐ��U���U�Hp\�V����A��$I��W҆!���P:��F �C*$��h�
��G�R$$%�X�O�}�zC�	�[%f�����������Ŋ�|8\�2��$1���;�~��u�3��:V4���f`cl\xn��N�͸x�3�H �Ф��Y�V]Z=��o߈E&�pH��7���y ���eeE��R�OUς�r�xB��Td��Po�eggojt�*�)�cґYaUSDyd�vr��w���ib�I�z'ݎ��QWߙ�D=₇���6�]�w���}�i�y���
Z�A�*������0 j����{�@M����d}\����������z�O���y�T��+<]���+�'���S��Ȁ�uA.r���'���8	��"^.�fN
�]L̖�@�g]���Z��hEH�n�O�K��	Ih1F_IIU�"o�z<����o���`d�ݻg�3��N�rB����ޑ�����r�.pڱ��L��x7h�d���EM��t�w8z�r���j;�w�\���.�A�y-}r���.���9_S�Bk��ܕՆ��,� 2��*2����ˣH�?5XK�M)��G�,�,d������s��n���Q�^~g��qZ��ϩb�����c\��5P~ϗ�������`TN�qd8�wHz��*,H~�_\|������������Н,W� F����m��ޘ-Չ�ٲ�*�����wSS�ͮ	�?�X�B���s�b=���e�&��Y+��{���rw�̘�M�XJʻ�l�)����QQ"����<�b�?����=<$c������; ~��u�������p��d��.��,���v���=+�5'��d
�V;��;����qk
٢�.M��HJF��2��Ks�B�m���geU�'3�D���)�1<�����_؈;�M���F�F�h�Ā��uw`R�E��<�d
*t :8�=6<�����-f~���s�|���eR�Jp�%���YVI����gC�|$� ���	��>}Jk@A?�<)����S��*�V�FGS׭H;�g0�,�����ѧ" ́�P���`�lG7 �@%��PR�|HSQU�Z���8�`Ć��=�_|y}T�ٱC�?y}��g&Ɣ�]\�y�9׳"i����&o��8OO��-�����խ*����{ߑ�������s��b����E�FX��iR�b:��BB,K~�MAG_ih��j��z�]����o�vuc|�_')y�5)E��zÉ-�Ro1�;�9���la�x�ڣ������9�����g�����l�9�@P�uL�| �Zf3G� ��Ȑ��111��Ƴ�-��M`�@���+��6d���l�YY{U~ϻ��e�˩*����H�m��
,��A򪾾�p\a�ͩ╕7t̸{�z:�ީ�gtSc�gw,)f���j`�Y��̌��(��U��|)��&>���SC@��0�/�BW�`��0���2�������S��R��U��x4��C;�n�R��SU��SY&Ņ��]���p\�ˑ@��6�T4|�Ϊ�73����0f6�������ͳ��&_�.�.���#��+�߇�C}PQ0	+���J�z��zLcԧ��R�qS	��s#�Y���ڕ�����B���ge%�)�,Á����4|�[`�B�����3���2�KX�� `��A�R	��ͯ/����zp:����g]�݌f�E��!��i�-��e���mL�I��?�?�-ཱ��'�K�z��H���U&q���Q��10 MOO�[�g�}g�3�+�.3t���p�ʒh"b�Ѩ�$�]Z�'�-�(��Wp�������s��}�����$**j�x:a{Պ��	��;���Ϯ�Z�*u�p���ග����gH@7}�[���̪:N��򇙰�sC$ʿ���5�9�.��L��^k}�^�!S!��{@#�&:��g�eN�����r,�(~x���z ��x�N6��	wI0wd@�w��1}�F��
4Hh̠�YZ�Egl�WEym�_�$L���a��Eq�2VN�H�r��s,���)
4<��� �A%�e'm�l|�����< f� !�Y�$��vɝ#]F���~�ܢEG�2D�j�{��`;����8 �y5r<(n��
�.Rg�M`��.�q�0�j`q��Ƞ�ҵ��~WM+����ٴٺ������S�w�&fk`?O5��%q	.�`��~n�2h����{?��7L(�^YXRUM�f�����q�@�.ㅇ���m�}~��7={�������֊�ٖ�ì�ۺ��m�`U�@�T��uZAKO>�Ż]�\:ɳX��a5_>���.�"e��Ӳ�� |薶",�J�ɺJ�qrC�[����'��=Yy�c�y�-�gĸ��O�R��O5���~�Bȵ"�x�������|�AM2{�g���'�u`}>LQ/##��WZ0p���Gs7DP���ڝ��/�~᷶�
P�K�8t2����>��)Er|��;�D�K������/����V01����j�.A*�|����IPW�m�1x���g�E�]_E%S,,1wo���Kc�9��Iq$�5����V��v۝�1���5�N�~�D��Q*�K{3H�2�-������_7���iɡ�o9��2$�������S�W�4����ϑv1���[)m�C�<ɄEy�����]$�a)𮤍f�md�~o�o'!�����u[��d1�g��}�3���� ]�z�8� �oʳ���D�et19L� /�9�s���l�E��ձQ{*�z�{%�;��� njw ��'����l󤷎��7Y������45r���b|�Y�����pힷGw],�Uq��S9s.?���T_��(4v���[�(���Q�֖ޝ�0װ[VVvt|\1)r��Wj�-�t�<�GL��q�z������@���(Uq�����h��FX��#)y�5iiI�f˳<��¼�x*b�4�����q�����7Z�	�㳲dd����kkk\����EBGB�N��_ ��o��������pڣw|�(u�ڽ�4����~�*$I�N8�I+l���^'RL�@S�.!&1����[nOh�ֵdA(z=����S�M��Q�Qw��S�E�ϷdTx'C$4%A�n�p:t�1��L����$�R��sua��rSqQME(�e��7�I*��oS#�8Y���Ъ�����Б�5���ԫ����ݺ�+b�LC��*㑜|s�~��?���^�Ƶ4�0I�5��?��~Y#I����h9�f�&�91��!O�c/yh�XO���ؐ��D�3�ݽs����̑��h|+[ii\�	�ͼ�4�M%�Q�eRa�a��V���R�x�j��jD`V���E��@9�1k��R��|QЉv��7׫�"��Eh9�Nt���&"_���nJ�_�(5;�� 5K��g��k������ִk=Ȼٚ%`O���h*G�� ��1Ow����ѝ��9�Եh���:أA��X5��`4'��<��1-`��輐$Ij�&�#�z�t���-(a���m�H�v�k�VR������TK5O"�?L�E�����s��Z�s@8vo
۠Yz
N��g=�L�����yx�=��> 
?iHΏ���-�8���]lc#��9�T
5%�U�zҿ�w�	>�-���U��^`��4LQ{ 2������y����������m�4�2I���G��{��㛆Չjeҧ1�������%,���#K�667C\C2�$ ��G�@�iW��"75�u����fFb���}���5,ӕ`CY�F �b��5��_�3���t�W#�_O�tkG�S����7,���ڎ及|z�h�J̒��L^������<B�p��D5Q)T*p3�/����N��J 6jg��]\2�:Im�!�u�ҵ�X�c��}= 28-<4@�啥�^��'�C� 
/㉒����*�J�%��}(���N��O(�c�+S��zD�a ��k���S
H/�3��O3�Ձ[��M���;��|���d�Μ���#ZX���S�~�G ���*��H�����Аљ��K�k|�Ԕ�1��$q�L�-�7���g�B�t֭��T�(B��\��#����!fY������셑���;�N������N��H {�N��)h�N�Q}"�&ǜĉ��/s� ]X�����y:�C-�����g0Y++ہ����p��d�اP/�SF���5ܶW���[tt��"��L���~d�]	�pȰ��(����cL��rX�gj��8�5�*�3��^.&	6�$�1��98�QPP�F�8!�`��yfO-���І ��%��٧���B�vF���K�j����߿=������h��,<.[�/=�Y�V���kL�޽�����z퇻��1��uى-���&�IY���2�T��5Y�����ڍ����E�]�`�:� �����ɉ�t&[�]6O�r%4�+o`a0�	��N��)��n��My1^ϰ�*��81/�r@<�n.�f�E9�	n�W@�g�pZ-���������WG�F��dE�yU�ˮ7���:��h�����&�w���)�(UW�B֕Qu�O��\Z����o��[ؘD����Ք\�;�g��<9�\�W�s��}9�UQ��߰��d]n���}p���~��k0Eptt,�&b����^���Ff��v�V��)�`��1fZ�b�Xf�hbH��<����=h�MZ�����i���x�Y����J�I�%w�qɇ=��,v���'޻�c�6��4���`+M/˫��������o?��� Q�ͮ�ߋz�'_x$�;����bdR<�xy	&RBc�b-��� #�L��F!U�ŋ��ܥv ��K�|zxT��-��nՉh�<�����カc0C^����z���u�pwq`��#o�����E#E���I�� �	����F�~�JI�X��Ō�,禅�wAB���{�X �����K�2��G��U�ގ��<s���c?��X�j����`�(��6T��^1��2���ڵ{r�����g�u��8�-��06���j?����ZxLKKk�z�eQ��#|d��@��Hyr�樁=b��Yoir4P�u �DQ�/ Љx�jIu�RsF�hܠ����?�H7���UJm���(��-=B�W�g$.��@I&'��2`�S���/A',,,a(��{�9$�X�U�����j�F���:x�|=7&[�_ش *Rd��f|��ߐ���b6kーDf����^n�8o��Ěh
lM���{?~\qK��<}���1!���]�	��0�Jn���7���>���YV�1�g�=�޼g��q����vO��A��.}ކ@��^�W�
	�9B�ݼ��V3D+��5^x�������A!o�K��r�ȁ���1�����8���,	+;;Z�ar ��5L.R~����u�E���B�����v* ����*i�� ��m�:U4��c����X���Xl򎀑n���q�3Y9�s�X��6�>�r=ƹ�uțN4�G�R���kjw�9�A���12��J� �YE���of��ee�?/�
��R���o��,E7 v�E��|������*s>A���U�2K�����\�?hR���;/�|a��l0͹������S�-I7x�2ڰ��rղc�w������1�!ݯ�b!S^fUX(Z�=y����%�֛T,&(88��v�1�O�"�9����u��X�7S�=E�F1�8��=�cD~�y���,�Q����q���S�f�,����{5�LG��^BV�M��ƜD��?Ϡ��$����
m]�֜$+7{�p�oa���:yxcb�cV(�S|`j�B/g��иϘ���yP|1�9�}`��/F�Q(�:��#'{W+%�TYٽ˃�Ž)�j�C[K��rE�
Fv�}��7��sO���3.�Q(>�=����)�`�aa�I)��v��w�9�'��1>X|y@(��Z�̕WV&D+��2b����|���L2��t�LK��QvMT���jß�x�z�s �|��x'�=��W�В�K�̈�&����Μ�S��t�'@-h�^A�і����KV�8�G���$%��.Mw�q�7m������53���h����Flw���Q�0��
?�������������r=���WP55�IS�?5a�����C��l��c=�Epi#s�;�y��g��v�b����-� �t�M��r�<8�����:4Š�r�eh1��m��B,��c���2S�TŃ���x�U��:\00����hXB�I�Cڡ6��B��X�u�S��]��= �5���{��%\�[t��<1"�>)?�#�y/w�z��@u�N��p4�sŚ�>0 =�f(�$�b���~�4�Ȯ��ll�z�c��Z��0dE�\���G`E�7@;d/��|6��8�D��
��(�����V�ʒ�XE��J�K0�_Y���t��ʴO��2��fEV�e�vr3s/�b�:�x��^��������xh�Y���QwU���;% �ʔ�ا)\�(��NO�u�i�����������`dd�����oW�RU�{L�Ȯ�Ƚ�Z�,���Su�+�5��<>O�����k��m�j}-mtq������3���?��Tk���t,�+hx���/NY_`��3�}:J<E��j��0|��o����
�_�6k@'���}��BL��ϑv2�fZ�+��CMVA��kN���Ђ�$7Z�.��M��x��8�]'��������^�U���^И��&�>:�.�Ʀj����������H��vI>z䍒����A�ԁ�����qv������$vE.�'�Eg�/�Hj�������ĥ��<uCK$$<,��'M�Sl�BX]��oi+8b�6����<8[;:�U�X�bo�ﺕ;��a����ͭ�
�ӥ+����n~���SL{�T���'�����`پ�)��Z����R�`E�CL�U��-yg ���{w�-U�C���0��F]rg��e��B/\N ��K"X��+�A�vOddP	U^����^B� �o��|a�����>b�fWW8�W�����j��k�m���;��y�����3{�v�J�GY�Uۂ�}@XYZ~ed��}Y(���a�Gͪ���_ع�Еn7�UD�,� .	5�������}��*�)��t���E7x�?�N�ߎ��Yv�e�yP��-�!~�½.k�Ƕf�RC�ZO�'0P؀9�%i�B5�'Z:�:�i�&����x�:՝��ݺ@�1��w.*�&��,OKC}�"_���1g�*T��?��nw�8��D�I��6d�m��<�Zxp� 1Sq�`��8OE�����9�0�G~�s��|1�OyU2�s�w�"�'e/�6(�o�������o����U��&��GG$������'V@�n��|�U��,	��{%�`��/R�����	��2ׂ�F�M,�B��09h���&1�;�m\L`Nq|�z��P��_S�h&��/�ś�-@��j�W��Li숈���{P�8�a/E__/5��~%�O5�ڕ�l:���vߴ١�xJ���795�wt��������`�4�o٫kjjju:�Y| �[�-�^���Q��v��]
p�L���G27@	�����W��ת�p� �y�����Ng�s�v}|88��O3��b��W�5��a)yQ��.�M#gﾄFy/O�����z
C6�\" !0цg������3 �7gg���1wo�Q;���v2��*�bL�D kQ���s~%k�'Yw�f��ơ��y�2��n����`k��P)Q�(�Y��f�����5^���ז�05?bȐ;A��(/)�5����o������=���mdRav�����=9sz���'!!T�.�?�2�/Q|��yav�kueeEM�-fs���z�H�M-�R���*.-o6ۊb���ʑ|׭i]���{w���s[L���zFl�_NK{�u��疷w7�׵ww�	����٢�767�ԭ�B`&��-3�Q��7/_���qPto_�J���6��ݽ�`"d����8�E�^�f�p~3n]k�.�ic=+6�5B���I歋Gq4׺f���[�OQGM>B
S���y�I!o�2W���EڲJ�Қ2J�` �bc��	8fP�ƅ�+Ќ���[bd��;���H̢/���5�b:>hE�q}	PF*_����>**.,�q3�D~8�T�V�U5U%�1��׻[#*驉m(�`�ޱ�n�!�����[m�q�YQM��KYu�EyeQ��{z���w�%թo���-�0i�i�4��mL
腖TI�-�hǥ�
\mUhW(1�&��¿��/G��R��+W,�!Is�+��_�T��l2��	&�3�w�^�˩7;ܐBP��`aa{�w�jı�z�zyMp�-R�n�':�i�㲆ݺkp��3QE�꬏����U���fr9��X�EC�JJ'�Z-�yuu��J9�x��Tt3���q�Z��hJ;޷��4�~�>�=�Sgt�gNd���Kk&T�k�Yg���H^m�'�o��]s'}mt
8�[X��ۯ�=t;�\���J�3���[u��~@p)M �$Z˿0��u�Y�J�p��b�Y3{J[��jK�m]t�d����.���.�֒��޾r1�g���k�c+%��-S��x�ۉ��}a)�W����r�+!��~=ӥ	!T�W4��c9<��	ƭ�B%]�Ot�K�3��%�u?��]4ON��m~m���QMGQ}񇣌��v���nH����Yg�].�v��bry�9 f�w-vN��M��d-$,\�^��׋����{���F���C��h~��~]��Ȑ��B 3�#
���477/쮿{��Q���.;��ed!��!����y&jAyt�G����S����/�?����o��$���??���$R�č��`ed��n��<����j��ӵ�V��	q.`Mz8�~�x>��}��CWo͜.�ڡN�q� ;���H�ƖR+D���f�8�J`"{������UXH�P�Ք���]Z���t���R�����`�X��{W^��f&eVς(�{$�kl���b�^�����T��F�`Yf�Ȉ�	�%Vt_����,�i�A�Z8wBJs��&6c#�I���^}�B߷~�`LR�*r{B��\��~H8Z�$$��|p�9�s;��ǰs��1�:�C�|��O��A��I�~qf��I��E�CX���d	��4����>�7���f��t��2���Qy{�������H19�M;��G��a�_����5*p��MR�@�Ob�_M^�Gt���5YR����5;����8]�G�-��;�-E�fu-�rQ��$^�a#lp�q&9;�o��j�Ո��?�		�t#rbWǬ	�,sf`���˔Bݱ�\z�]�3��gI��	����%���2��mO��|���x 7+��D�^�ZXn�1cfP��8u�_#��@��u3s���v��;���''	)�J��PY�ly�f�͌���G�d���<���#���"[#����t�ej�'6���{�~T��b�+�M�&815u�}�N6R�vPj	�"�P��Tٙ��I<RRR����N����`�����#[Ñ�c8��,b{�W~?��$)��,{�A����������41�����.��D�[s������'�����u")&�,�9��!�@;��,���MJ�^�����6�݁�O��/�7�:�5��0��������(��5�6�p��< �۶p��������ƖF��ϋR���_�7b�@�b��zV�Փ3�1��,�˃4��T�|f��!���H�P�ASr�uP�������Ђ����Ź�^������Є��ɡ�A6+�p����ǔ�6�U����Stz�rK(�9ݙ�������U80�Xj���P�b��֨�����p��_a��8�:K�_?C�,�$�&�~cln|�,�x�N�m�ǒr�]i���'==�<d|ĺ�e0����t��\m�d�V��@��v]O��[[�����@MR�N|��$�8��1D��^e__�,<:�"��
�崤H�ЧF�M��s��j���j
 �z��! Q�� ̮�)��j )���v�2h��pb�;9=���L���CL�g��:�1j�@�8��wz��ى��C3�����0��b��!3��^vs���!�hi�l�+3���}|�����������0�]8��n�
�Q�g��g��?�_!��u��%���i���䓜�Z6���DF`g[n /X�3�ݔ&bzN�ċC<��E�EIM2��/#3���o|��q��24���ҧ:e��c��݇^Xt׵�@� �[k��=��JSq.\�4Ϸ��o(�(Y�����@(2B�WQQ0������Z��wy%��LL��E���1员��A[Q�zm0\(��BIWU+��Z�РEDa�ubne[Qc�kh8�BA�ԧ�;<���T�l�L�N�L�n	�?bD>A����3L��Nd�����_�Օ�_~k���,P��#	�ݴ!��������0��,?}����!�ɀ����񐜒��h��H���ɶm{�7�m��6ۛ�͵��l�fksM����{�6���9�s�/���fv�y���6DpVim��~p�i�onx׻7a��3�T��F�jG�A�s��\i�^�^F*3֌����t��7Ӵ�2.�2�dؿ2�8��o�ib��R���԰x~�ψ��J �5�T���"��W�]���D�n�& �TO"5��,�z�����L�s㾎��~L
2nl�z���	��L$����w�1y�+�v�E8�Q�ug�W5<"�S���?�I�u��FF���O�w0��;��� 91U;,,M.��7����!���J�Aڀ$�����!�$�D�-�/�#�*\�O�D���m��&'���n�T�'g1���~p��Z�2�tQ
���x~�O�/���S�+���p��-������xF���tr����D����t�dok/zB͇72�QS]�h����{�8z�o����u��wӜ�wx�vc�]V�}�^���J�!>�����1<`����;\+�7Ű����TO����;��vcL����&Ҝ��.��aI�s���'m��:���q�/+uR ��(ܽ�W�ݶ�j��㊕�I�c���;�#cu�����ƀ4J�����b���m�Z{v����T�}����Yw�Q��yM���;�X�qH7��wi[�|� I����M 	<v�O�����=*�\*?�ؚ����0!��e��:�C�j'(3&�#=یL��A�u��6�Q�j����o4q^x ��X�$�.	�^ʥ�t=r��ͧ1k[��EhW�vkS��*l2޺�)y���KXa��-b�aw��:~0�ݶlհh���e���~dPip��A rssC�7;�5-\��db�&�c2M��_�A����^_�T���=��_%/���z6D2���@c.ƌ��=J������u|�wM�M�$�ёC�$�۝KDMu�z8T^V��j��"!#���L�~l5X�p�/�����^��_}��V���z�_�<?q{v?T��<��X,���)Ѕ	��c�µzK��LbԅE���vZ��1�d��5��*�a�����h~��*�W2 �$�]K��$<+r$}�ذ765�t㇋\i�_�]|�/�Z��^�9��?D9��ʛU%YרS0f�H�ؽ�0t�*����mDI��;���"~/{�܅K��)Ͻ&l/�)Xу������**����4SC��aӘ��~Qq1�g�ۃ�y�ƂΊ��i`wK�xį3)g��I6��я|�Tu?n,�UT���b�D�/�,��M��.,,$_O��T��Ԣv���` �n:WPL,���=��I�'
�̫ǲt}P�TVJZ�w��.�1+�u<�ӋI�狃�o)��<l��rR�X�[za�h�n.��\�x�*%0#RI� ����Co=2�� �l#��.�u�c~����>��CPj�uC_�d�NKE�D�n����Y_�Eb�7Ő���OR�x����)j���ᕾڍ�����r�����k�FA����O[����
�;:W��.H�D�R�`������:[����Ait��rM��$񀛳���Hȧ��3y��ׁuFӡ���O{2��2v�#��&ֱ����l���u�ݏ����5md�/D�p�1��P:�[���i�|�P�PQ8o1�/9�9��%�4��cb�f�w/E,�s���?��ݶ>.�;�o������C^˥cu)�뫴pG~���8a�6�F%y��x�N
:47�o��d�	'L�du��M��D�>mnn"�#ݽB����7C�)Cz��fM�(!����k��aAR�e�啩!�;EXY�@����9B>���F�r�R���:���m�s��8[�\��^@�x�.�q&<�L�/`Sҵb眚S��AT3������2�R�b������1��˔���g���t�P��?|%���¿�{�oJjt��a���8m	�ۮ������o��Q�p���/������Jۉ��o�о8{Bq��ܖ�x��Q�4��$�q��;��$�����FX�{�4�W�x��w�f1�~�un��f��;��Qtp��C���1�?3�v�%���E>��绤h�R3l�cVa��%}` ���P�ڹ�e�q�_���Q�L�)�uD���䭥&�$���ނpE���:,5���v�2��>��G��b�,���ވQ������u�8��ڭ��S8��n�2i�$��#��2qV��+�J,�샓s�$��I��Γ�tm7��}�s������x�����Dh���)c���	�$�3kJ�i�(���F�նM�eeX	3�H�p�/��vu��oU����z؉Y�ٺ��P�Mt��|�G��.��7��B��W��!�=���<�n~h�La*��<08FF�p¤��k����������͖K{o��	�D�M+z�
,[}���$:$��cl�\:/�������!��n)W{�/��e��"N8�_�K�������ד�G,ZO飼����q�9�l(�~oṽ�QRB1׵�>��O�b�������p����+��=���]u�A�a��>�O����i�e/arM�b���]Bx�b���0ve]/"��9r����m� ���EE�U��:�br2�<aD��wHY|׳�3#՝�����};=/�&���Uo�mS�+�s7Z�J��ҡ؏pNwq/z�����vM��/��cB���zf��pw��]�yK"��`�h��(/��3�����+�.e���U��p����_���,D����T��V��BR�HR����ft�T�tz$���21伃Q����;����F���%��}��q���4h�^sgF슆��D&*�~Zd��׬����E/�q��8�(Ϊ�����s�0�M�Xn���ʴxjW�rX8��b0jzz�>u�ǥZH}{��4G&z��:2�Y��8�Y�X8yR�=-�q�*�za��S��aKZF�9�6bb�0�3�ՙ[�˗��r��<�'$�4?װD@]Q�$���+m�f�y
��I(�����=������s�jQ��'��s�iI��!a�XY�cgG��PہL�	=%I��lDp�;����*暄�N�/�g���s\2�mrֲ�����ߒi����B�R&�����u�Ѓ�6�����7dLD1�W4oTi1{�#�i�������?��F3;P�c̋���3Ɯ�fe��G=$d���ka��}\s/§����=���
���� �����O������_�:�O�CD���G��g�@�o����?G�ի�n%��9~��F^�{վ��g�455�u�������
 �8[�ǚ�}�KS1������n�(�py�����D���9��"��d������&P�.,���[;���=����a�B\`������1�H��-���6\^p<l���Pl�PN��6����<�2Lt�̀s��Rl�� .��?9P�=;4�{=H/*UF��bX�����[�iB�Q��5�<�p�Y����:���odRQ���\]��;����#�y�>x6�<nߢP�M���r�����W+� ϗ���Ck	�����D���k��o[{ά�<Q��������g�,�9��P$�a�*a  e���|�Y&� ����5_�����Ԑǘ��lkkg���]'���#;7j���_^�M�������Dg�'5Ģ�@?%RX`��w�6� \8�ѭ�����<��o�4W(B�W�g�$PN�4EV�ni��[S�g3�$ m;=����?H	�[L��fps�M,ʦqp ,��W�\Mjߕ�����(�D�~���a�?���.��^Ł����Ἣc?\B!5���}z!뷱!��<9��7����Y �$5���pm=�6�f�b�0pǱ�����u�׺0��+sF��/%�][��]y��Q�V�� �y��#x�!����	{l��$����v���5��e 5{[Hrw�|I�7�.�X��*.*o8���z-�E��pJ��Q�9�JBزs�ZԞ���Q��0O���[��mvm@�^2��A�a��Qxi��ns���b`�XY>�(5g�yި����G����X_����T)���Ȱ������6�>#ڷ
v��@K����^�;�����}�*�����7�-Au3����k�ӧE*Zi~���#c�*5S�7]:��+X�,Y�S����V���!ծ��wVr=xQ�6�
K���>��B�Z��^�N5:�������.`m�qBd�vl��c=�K�ҵ�"�u(�w�d^-��*�����=0Zr}�Mq�}�Ӂ9#������r�Qd����{���wtT�rHt8n|Qi�b�S�8�:^�XEb��m�e��>\wVƥ�Zޡi���m����zb*��I?�y��Ӭ�J8gxE�ޘ��sj�7�תmH����Yِ�����.l|xc�����Վ7��i���uU�j8��z��%J���O���u_�|y�
_�&�VZ��vK�9��~ )��}r�����_q+`$ �)\���* N?>mø���Y�SW�[���A��>�k�9f`�oz�;C�G%&V��H����� ~[�qHkNNF��zP7]V�|<���P����P��մ^^V�p{��(�=��������GJwxSڤ�0�
Q���h�<�|^ף埭�ޝzׇ�*#Y����N�u��<(8تem��j���T��T�Ү���5Q�T�a��?ǂ��~���^0$��$���Q�D'R�]�H��R��'V�ʮPE"�\4,��
�zp���jѯN�_�� �A-��@�(��J#�&���1-]Y�����3��� �����b��ݯ��2�!mp|1��S��������k��)h�*�v9O����i� ����R7op�MV�5�aM��d�p]E�z�K�O	p� Q]�����h������m[0󮲒��|3�����E��0��?��µ�h��J�u���G�=���1#G�g�R=��}t��Vc�`A���zq���%*6J-�Uŕ��JxF���/�O<�t��<�.�-�����%�C9>�݆'F�z���q^;۳�hɋ�hZ��5��΅/��G���� ʃ���F�|�U-b>��풞E�6Z0�fc?�"W����&PaL��5wQ�VU	���3Y%4[����h����:�$�#���+��(��i�X��˿��i@�$l����р�(Z8�h��(�C�lQ��LhO�7���B�X��ȷy�%@͆>� ���p~���}������!�R/5ɸ�e�;<��x���Al�;y��C���ƿ���X�YV����츅�1!77E��	W���e0�i!5�ZdU�V��k:�M�wݫ�F�$������̶��RY�L)�{�4����׎�Ρj��T̽HD�'�=��5�R�aQ�{i9�\���` ��Y�����C�����d9`����Р,���L������ѧ ҆�ψc��b�`�DNW��9%}�|9����h%W�'��6M㶪}���� �A �U
�W��ʓ�6��z�2���-�gҍ9��V
��-��tc���B�C�c4����B:4��"��(B'nHw��Cs	�1O�u_!�5�F�h��6��p��7i���~%��f��)2H)q��%�7F�۬����9�)���(�C<H�����f$(��ymXec��)ab�޲J}��e54��du#��aa7L~KS&8ǟ:̩/;c��|J�s8ftyw�T���G�M�Aa0�v|H���3F�G1w�d�=T���V�|Lo�qp7G*~d�Q�|�B`�4~�X�r����t�
��
β�f:�9Ǿ4�%S����ɫ����o+evֵ�u�e�aU/�)m@�a�	IW�0}%�.�!o	n;��m��c�s̕/J��2I��A/]�8/a�Ы�
��ox�ܙQ���DTV��`N�	��t+�� ����ȫx��I�Z��0V���=�}`"w3���$=�l,J�>d�ss���'5Q) �9t|I�%}�+.���r�1m&����'��
HnkfrFЦ�<���p�,�D #eAy�=��?j��!wR��Q�
�����~�/��Vo[X#7����]�6�p��(4W
S\I�]Q�'2�! P��?�x_a�7�$5�$�h~��*5�A���E>��vf#80p�RC.*�7"T��.<�^���ת�G�j�M�S�!����]�[9�����X4��$�
���a=h5s�,�X�1I�U㌁�����wR�;�_LK�f�f�AԂ��8�G�¬"hذ@ܛ����]�F��{(y�s&�.kǰjJI�u��YQ�d
Ŷ�F�{���c"n���'����ވкR
Q�B8!@�˅(�>�X��,�7�bC�{����\������H�s<�'�o'�c�֋��/�ʤ�U�kR�b�P�7NQ�c��1Ș��{!�1�Xi@'#++k����b�[n�v'��-����i�,<��G��$�t�i�Fs�[���VX�p����Z-�[~$�1D��2�hNx@!	�#�b����c]���W*/[�;T�vmn��RP��z�U/�Z9�e����5����9 jy{Y���ιV�VP��z�mV_�Ŭ��p�(b�&�:6��<  0Jz;brM`%H|B�Ӹ�7X�Ė�W���+������jMr:�ƨ��H�X�5��ȓ��c����.�1�����"���N�X�)'wu��[[>s5��0�[GN�-�/ʃG�@l���K��L�)f�
O�����T>w�1� �xL,0�~k��T+�UG��)T�~�~��5;F��f�?j��}�� ·ҤY�T�ɘ���A�:�Yf�<s�1��	��ί0|8�U͗�X�+p���
{$�yHq��ڽ��V[�]��}^�^�����/�<)u��m�?p�?n�c<��wI"Cl�N������쉅Y�e	��gP�l'���ɩ�ߤ�CE�hA���c!us���cv�&&L�>�E.�e���n_o�؎a�p;���_dk��b�{�@�-j$�C
od���p�s�鵑��ھ*8� ˻�O5���A{�@�� ü��7��d��ʻ�U���o�>`�ǐ�H� ��I�k:���W�p��wEl1��u&en�X����y���m�W#ҟ���B$�F�6�0��5
�R��s�䦠�������>��ۛD$�}�Zwوp7���誒X:#�W`�b�)/�.~k0eUԪ� ����x�ÿܟci�Z�VѢ� �4�
r��/-ݽ=�蘒�I|J�F\ޯ	���ꁖ�X�o���8W�?1d�t�I�v��OFv�o�O)d�o����
�p���w���J���1���a�(m���&H9n�F��A���:xV�Hp��/f��\�D�6C|v%�C��A��?��%�Α�^(��cE������"��+\����<�IqEm<6��XM��ʣ�O�C�Fż�S��M��L�0A���U l����L��-�S�i��6�v��p�>����D�Q�u�~�����eq��D�՟πze�����At���A(�Y3��L@��o\Z2�����y=�
��7!a�·�Y�26x����I���2�\����Ed�?>/p��*.9f���|���3I(c�j���,N�RE���vY����@>��N�#"}���p�e#�� �f��Aq�-��|s��iq�"��a� tV���C�5��s$:��F�h���*8�b-:����b`�J>1_(XsUi���K��� �Q�k�78�Q����R����j��x����Q���n�6�~�`��ǆ��%���W�t�t�o�d��t�U����rs�Ƅ�m-0P�[Jh{��?�_�3���{�jЪ[�5�,���QFh��sѥ���Ӵ�Aдơ5�(<m��.��z��J���..���c=��=|s����/�+r����9��������'`�7�Ɗ{��nlĮ�����]���ڪ������\�70�E@[�;I	DI+�b ��咱G�c\��zv����$���_4�D�m�t�(B�m��u�h�bz ��I�m�t���e�79K�(��9����4�Ӹ����GG�����Ola�>1
�N�|�ܱ�y���U��x��hu�_$����0߫�������֩���GB4��U���z�Wiv/���[c�������S��F������#�ƿq`CZ�[z}�q �+b�e4��{�Cu #���D�y�߂��Y�H�B�r�ц�J����~=8H��V��xϷ��t��Ђ���J[�@�b����Hl��28Pˍ�R�����|���[�F�H�ۚ�:c&����s$Z�MW��#���n���р!>T6�Sa��뇗�d������K�ǌL֋>;������E�M����9^�Ҁ��do���2�R1�p�a�;���QzHx�;r?��Wu��WzN!�:�~f�/�`NF��8Ąr���reOB/���?1UZ�5�J}O��e+�K����Q�!�߾9�⪳~��CʏA6�6I'31%_2Z6�{&{��H�xt��^�G��� ��s�-&����� @� T>�,u�9*,�L�>�8��+�	����H"�������6��Ʈ3�&��'��:{����'r ����.|`^^G[ҡ������, ȣ��&ZSE��+�me�q�<|��/\����:���5N�J֞�Js@@�Cv:	�?� +mABh�&qP���5��&�*��k7(�E<�y���[��B&~��MD@(��sH�`��V��#X�q�=	�Z}ƨ�J69v9"d��[��m�G&		*R|��OF
��i�%:�ou� ����� 0�X���`���d�#���q�19�sD��-ڡ���!u�Y�Y�`�kS,�����>�;��?a6�to�i]����������ɂ�ED1Q��m#66�k�����\V��vP~��<!�W9�(,y��/ �.�f@`�[��~�ך'��MG�_܈a��=���X$>�X#���ƚ�8�)�?�%MRV;�_�*�_b�:���!��y.Q�S������1ND/T����ڌ�-�����jC��d5���F�	����5����}!	�Mщ��>%꺳��ܡ1^�������A�Y~��X|�vˬ�������.���ǯ�I�8%��S۶Rjz��ڵ�%�I�A��H�m_��ꂂ�ɢ�E+��3��Q�ݑ�^�JX> ��n-D��*�l����~'cֈ�;�9�<��ﺢ\dB�.{���o����~�͍
�IԷɟl"��.����)�F�U-AJk��s����������O>�q���}��޽{�2��j�ZӴ\��P�'�<���z�$�`���������]�y���Ž�H=n��Ǯ?���?'$�`$47s�=xa�/�Z2���Ȏ9��T��Ӛ�����$��*�h�ɍ�J��`���c�2~xCJ&��u�⸳���q%��Y ��߉����#$�b�ǥW�;*���6ւ�x:���/$�m��1~���B���+J��d<q�"'6S}�������\ꁍЛ��qŉ��IIc�SA\4f�!	��A��>r�ش�*������.����W:�!��T��k|���)��ʦ���N�V�t��wR�()�N5�<�A|0�h0��s���eC���S����C����*:,du����#jr�L�y2��m���g�c]�??�}��F���y��\�\tX�����p	'�
��,,qoje�cܨhuf�4�kVgs�:���Y#΂���SyB��i�|b�܃���ֻy�f�եf�����pyJ>.N�|�kUA�C/-x�T���2�;��( �4T*��Ѡ��Mǘ����C/���t�4 � M�G���E���q$\T:�쨼��gN%���&�����CM��F�9�d^�R����9k#������#f�¾��9�<��1�������noD+KR���!�a^�`"���]��'��|���rrlCig�K_��|v�)02���}�
7 5;q�ݝ��]�Ɔ;Q�>�l}7��[�iBn�R�+E�O�gY+��������̰PE����U�p�0:�q����6v1KҺg�X�{���i�=���Fsx�E���� �V�/����@�VH�cOĩ���������;[�A��VUCTj�Y���i
�t�����Inv������$(���=���FP��K	N���:̆���ԛ�Ë���3��9�_.�����������,�p@S3++�y������#����j2�8��nOa�p�JR4�7{y"}`�?��m��h�踔p�0j�[�@&��5�b�p��A��'���lA�hﱢ۠����@���{wr��$v,N�<�ә6�<�9jKe-"*�0	�	8m+�1����Tx�}����:+	O�Ձ2�h?QEŲ?�u��3pv�����GϟZA:���3�@�5����5n/qv�-����;}[���l�gl"=��aa�:2��A�-�f-����J�?�{>�8w��������4&b��^���I�����:-�����VW�TO�Pw =�/%�������<v�DYq�!G�x�������l\�Z�=�0a337Wi^����55R����ou_�4�����������C��9� @�UX��^ Ƶx:{� ���y���	�%9�Qq����t���V�P_sۏ4��=�j���#Hօ9	6��(%�覧H~G��ݱ�3&� tnB~�,��N�a=���pe8C8#��v�:�.GAaf�PĖ'gǬg#.��{��jjs`x��d����f��O��=vVg���XNi��D�KN�G?1��>�ĎR�}����� fZTߎ�(ɞ��|���xT@�����mKs��_
� /�|�q((�Na�a`��n���+���F�ͻ��¿��
>TO���K�����l��|x?��Fu�|[[)������� H�=��3�QS��9}'8�C�-ĩ�i�������+�F-����X0��z�El̐�����"Ŝ�fMr8�5������Or?��#{0������tg	g�9o�2x9O��I��!�c�!�O�l/ƺq&��Z�sS�H��K����lCsYDc1k�R�8�i�]���8��〡Ti�'4��]�� �0���f�,���)���L��o�yl�L �<l�+��%�i�ddd��w�����y���aSR|���يۃ�R��oW�E���b�,���!4���}.�d�\��nDXh��/�X��Y�6�[�3�C�R�����&��C�[k��z14�\h��cC�9P�S�>3��z@LY!3^��3��F�V@6�}dxbN�K��7<<�L��p_�u�^���4�[r�-����^�zĉ���Y�V���:���f�k��$�C�tw�t��L��h$d�km��ȟvW�*6o��Ax�����ȓ�G�$K���!-����/��̟����ËH��م����-^�M���|�~ǁ0�-|�O�}b�����כ��k1�	���-�UZESF�0���� ��]����$yh��l/4�J��Z��'8�H&�P��|_+���roʏ��#�}��q�d���R�w�	YXa�.\��yZE/�����n�q6K����:	J1�Z�,.�pb����/�,V��e��h��r��7�I��WBP��B��/d'=������rr����w�H%W2�o~�AI#YH�UUmM�K��[��!/@�r0���$Eܺ!�R�W��8����ă[�D��7E_�s�����;�U���
f�:�sa��󟔇]� �7ֺ5"�<@G���vd+����A:K�-6���5+Z�t����\l��ǥmM8M�t�iz��T\���wJ�~'�Ժ{�Ҟ�G�R ��&�I��Ke07�������|�^%�ᆦ-:y��s>i�f�HqY!&�NA�H��2Ū-
B��/K�iP[b aTr�}C��8�����Aq$����)Q��ѲĭE�t��b�D��������2��qC�Dn�+J�a���/��\��
B�e���y�+��_��hTec�*3�9�uM%m*	ז6�k�Q�m�	���'�tv�ëa��܅�u�����.���;�de�Y�(��x�E<^���"b��oc�&_�T�T��W��JIt5�<4�:�A�I !"ڨ�ƛl��	}��3)�U�bf������Xj2�P�U�%l������W��C�q�KO {����|�x,�SX�� Bnf�p�^�����(ҟ�o��ˤ�"�$������	�������������s�R6Z��!rY���;����	UUկY��/�얱�\D:k/G���pW��;��^�7*j� ��K!B��:�A(��Gh"W0����	��f3����ށ�0��0���ƿ�}�h���w��I��X�w���ݟ�J^:v��t����������)|ff�󊮺q�zǯ䞟� 3��:M�����Dw�����*E�j���
��C����8�6�H�����$=�aO�8��G�R�@UR�w�����i[��q������n�V�A6d�}�}`\ ��tq���=f�Bn���!QΛӾB3���r6d,@!+�n���� T�є�eޝ��f�X���tF�lp�u�;P��^)R�2�!��؎��A�
���y��OOO���������Z��GI��sg�?n�:��Qa!�t)��|���:�����M)X��Y����qH�Z�� x��#uP�D����5��>�GA��W�8���Ta�3�+���&9I@vl���%���aO���.{ I�5=&s������]�Y�7k]�^ޣY9�r8�	yW���=˩�����4�N�����KS�� ��Ga?��绿"��Q�-S!��}���`�ȋ^R�56o�x���/��2��_�(����	�1�F�&�cOf�:�SȡTer��_��,���^�5-�:1��9��^�J�D��M�FB%Ca��L��N'�	Z8Ek��&a��f5/��",��?uT,�C^������ԝq�A�������>B��W�F�Gf��7�:%ۭ��9B�	}/)gE�9�?x���!q�` q�br`r�eY�����B5׸5�����ƹ�;��[�Y��XJn~�b���1�}oVAHm <`N鿭�,"3�s�X��%4�q��ޝŽ)i�*�;4Ҥ)CV��/��
�����5A� ���>�������}�N��+���J~F�$ڭ8G-���al4;�
�?W,0N�ݷ�<M,�k{��J$!�P3D.�l�2��R�ǈ����2P0�7�b��zz���>΁�l��8y��}��:*���ȵ����)N�o(U����'O�c�[���P��]�°�(��T^C!/S�+y ����I�>4y�t��&]]�W4cU�� ��Ǖ���l�����b��|��	��l����\�ï��k��Y��.5]j�p� ��
��	�-���C_���o��,�Wh��3Y�=�I����?�F��/..��C`Qn���#M7v�\\��~�c԰(n�
-�'�����a��o#-1�ΔÁM�7��Zh��K/���!(�@%�=s �y��%����T�ͮ*G�77�:����R��l5f��T��J�����3'�⾉=-�K���ӕЪ�֕_D�+b<�ٙ��6j���=ɪ�͔���ĔNL������pCa1
���p�̑��+(Ê�$��KK�z��6>�.&�
އ=�k�rq����_c��ς��d��������"�L�Q'����𲻐J�*�Gp��,�W1�K�h~qXvߦ�£=�`��Ae�a`K���x?t�r�i�8v��̒��f��R�n$8j�Jz�Nʸ�x.rw�_'&��ƚabb�b$O	�Ӽ2
)2�3c"��t�ԯ9�:!	z���Q�}<������LM���9�}|�<�;k�?�W��璘j�-ٙQ�+£�Y$Gnդ��uG�o_�ߍ�qS`��{��������%-%��0`Y���]�)���R��̖�u�B�U˩Z���ʼ��|?�$��}$Vt*��@��4P���u5���l���E�W]���#|�b6^�EM@��xl�v�o3+/}J��o�[8ঀ�]�Y�牮m�,���ӧ��{T�صq���(�t�u9/��c�-E�=���D���z�,mvaU�����v+��5wA�3��V����P���%&��)�~X��y˾@��8�0-P�>�4�_A�Y=)���R���q�p/�?
ܶY��������b�c)1aI�d�!��.Ia||���w5v[�����5����$8���T�"��^_ �K{�6�p	��F+;Y��7J[��!�����)�t�@��%{��J��XY�պ>���g������.�Y��l�*�� ��<Ut��nh��PKa"�^
>���Z��|Mw��~R?v�3�f�6�΢	+)�� &���P<U��o�<�e|�?4��!��%/��z���K���a��j��nS#i���Y\�Z�Ƙ��9".��g�pb.~:���"H��6]���e�y|�9�{7�"�~������!F)�U�{;%�|?w4L���a��#�+TQ�ؿ�;O�0h���t�O������3��������X~=x `)�!	s��^x�����X]6��W��)n���{����4�W)���\T�|�r8��|���m�@3�@�eD�UQ�ʌ�z�=h�����5P��+�WϚ5sj�Ly��ʫ����n*6���(j	Tt(;U����x�����(錈�m�m7��S����G]���=52��VG�"���d&Ȁ��C>���0�!��Y�M��c������ύ�Ov�;���#��¥��vɠ�������BGZw����c�`�5��;���U5�Wy�����R�Q��2��^�WQ�vU�G
�\h��8i-�����AES�	�<�Ҍ�H	�1!J�ш?�/5�}�%��������@؎|���4�sW]m=+֭�V�"*%Ɲ� �9�~�\1��u��~ Ve���
��B��k1f�%D���%���e̪��3��p��	�l�>�����j��N*�-��!���j/;DX����kx�ѩډڴj�bם:�o����~�|�_s�#&Ƥ��C���y�E���t\��#!P~�^=�xl�dpB%��`�ؒ�'�=�1���fPGX��N5j��z�oZ�:re��������4��޶�HR�(aF���'�F���]9����5�*������!�g����\��>(fq!a�C!"��)/,�#I��8�K̡ �ar������;��9��Kս2��h"U�}��?q���Ʋ}�:2��I��ݱ����@P�]�[B���ú��nϫ�W9p1�a��i<\ re�;��A�Vk�R�'�����ߵ��{�|3-����
�J׽��slHO��6f⴯;�/�겍�a[��	�����K,��H��vX�ϑ=��ω	P��=a&r�oY�djd!X����->���ä���P�yg�R���Ҍ皓�Q�a�m�h��8�����{��U�[zъ{�1fK1g�}|)[��3܀���_p �������R��x�w�~[ܿ+%և����a��
�-�_ߙ�~���ј�'�zV�Ws=T�_�T��=�����k�9��� �����vqYa�5E�^� ��e,q�H*����$%AX[[3�x����l��掉|��ӳ<�ɯz���#����^;�7a1�:[2��#���q��1R]���F~4,T���Xм��!S�z�@�,#.��[h~�8�A�g��h��~E������^�wQ�T/�o��;=hL9��@,0�f�ݪ��%Xc���7%��&�?�/'g��1�I���9�$�-vě��8q/�����_�Q��Jk�Jm6H���R��6���@�ӛ#y�v��&��>%��W��H�ঞ~vL�*����2��xo˚����TA�ɉ�Q�1�����a��1/|m�+N�2EX����!��t�	6���Gf\[�]sߐ�C���nMo��)�̬�-�u^iy1��9��neȞ��^T�p7�Nk[Y�g�PA� z�z�_��`��X����/Y[�{��8m��Ә��c��Br�?y8�|ٕ�U��Ϳ�Y7�Gݥ:8�e�i1:�-��!G�QN����W{{���F��w�ɛV8���>��6�]�Pjp��_,�������}���� *���֦O|]�����)�\��{���+�*LO���b����(�>'f��&���:˨�ַ�t�t7
�)� ��Hצ��CB����K��A���]���y^���X�q]s������"9�-����Q*o�8���pDbn/��X���7�WJ���/���(�$�`|�_��V-(��n�d<P����	��z7vݦUx�h3O��s�8�b՞:�]����`�2V��xZ��&�\��&�x7�,;U1����և�i�����z�� ÷��=k�A��r�h���)��g5Υ���y���%�N(64$���u��T�S�r���l��հ���o��\up����ܙv<�.��X<�܏ڍ�u�d���P�ʿ��亿��q��S!-%��T@u,��\3����ZQ�L��H�
�@�=��Q�c�m���G�yS��m?��vm|v���X��v`t�'������Փ���>�f�l��Y����'Lc��Qj�G�Dl�Jq�ؾ���hmm�l��~�R�"�`~ =� �T���kvx����k�Ǖ��N��O����q[�cA��e\�r��	�l,?��<oXv���{�� #����5`'���J�i{vLd�X1m �/��o�@n�C�$#�kdsqH� t����x3�ّj-�J���V�K�i��-+��: >�0b���.ԫ�
��| [������ԟ^��>:�,(P��Gx��!~P#�)l$u�p'

������݆_�J�XrI�)��=�kU�n�i��Y�ZX�\~����3h��Ԑ�ʗe��Ŭ�?���ųqA!Yτ*�����j��2�s��i���C�u#DFy�ˊ��8�t�����OF�4r���q��߷ܮ��D܎�V!'���,H����@z�ӷ�T{E��ź*�vob�7�磗5CN8u��g;º�-r������\�x�y*IȄ��$�w� �H~S��GҀ�4t��Q���XXU�"���y� /D{ i$���ˇ�����ٱko�R�^��&,
ba����}��K�Y�B��k\:Qt�?�?�/ϳ�lo_+�^$�݂vK�����n�n���Ď}r�oNK��9~B�ύ�r��$�2�J``T�>���K�s��i�͈]������ڪ�B��B�H4ӣ&�~�o$1��\�о��b���'��=�m�+�^N!�PpЃ��?��_[{&��z�A���������g�#f�b����:H�y?���$v���B0�I�_�e��3q&
}t���A붶�G���m�]ik�P��b�v�1%>�)����yԈ�
:�I�9���?��7heaӬ�nMz����������l�.B��i/�ku�)7!�BE�*����U"������H��iߘi�����rKc�tNUUlM;����؋KřzP����1tU1w���O#FW�*�[���ϝ�����r��p�1�� z�T`u�k�웼�U��]�;��~Rn�s���.�D�����h���C�������J����߽����5��X,����p^x��'G�D���� e�0˛/@�=�s��LNgR��AJL�Y+�iD�~�������IA�����`�7"P���8�b"�W^���S1��t�L���6�ݠ����=H�zr��L��+�����$[��0'T�6�r2F�W��Q�i�M��t������NCCE�ʶjl@aRH)����g�>��N���
P_(�k ����E�/\O������J�`:&�V!~�ּ�GPWx�ju�P��6i��_+�u@/��{��P�����=�d۱]>㗟>��d�9�� (�UZ�.�Qqnޭ��mu8������+<<�t����¸2)�m��;��K �_�u��WS��Opu��q>�84�ktS/ <A���<!H��Đ�CԊ#���-V��o�>=~b�<v�#�E3h��:(49�[�`XX�9?������w�|����{nOV�"	�Qh�w�2Os��;s��7����L�aJ邒	.@ݙ����ANQ`���ByB3����6�ٜet��6C��Ztq2,Ժ������}�v�E��e}+�8ϩ&�aa��m`���w��홋���N�eV*��CEc3{�2���q��h�E��"h�p\����\���u	��u(����dqss����4�Q���c��q����G���w^P��e������9A�ߦ�tr�����9��^�g@���L���O��\]�M�M��O�E�킠���p[h6i�B����(m��!M�����&=�������_�;a �{����o��Kt���076��ؾF�55D�У�u�70�2q#�����a˦���Ə5?� �������:#J�>mu���cd{�ɀK���P�M�N�-g��}�y�9�P���Giie�	�Q����p":)���c�:t�_gd[�?_i^/ic�2�!�d����|b����Vz-��˹��
�1�]�j�RHj�RF��fV�,Q��Zvf&
�>85�ǩ�R�����?��~I� �i%m�����(��b��zU�}1��gZ����Ֆ������9]����mc�4�m&����\�Pn^))]i:9-/�H~�,Z�+*�"d��V�.�d�7���ܻ@+⨉/�]o�g<��!��YŃ��|�Q\p^�.%e�����ݥ7��4h����U��kT]�PöM��S���d�������p��$�;Cѥ���HĎ5L쵑�o�|knks*rss>[Ʉ]k�F�Z�5���fT^yں�9�,�+?V�8]b6�@6�p�c��u	{�{��&sN��ā��ۧ��
G&����z}���?���
�"�j�#GSSSU;����p�/'�����.�=o�WB	h��5T���l��p�w@��lz���dg�� ����6�tT^��Y��mM�[��-ui0>>!U�AP��n����2Qz�vB p��j�J�<�^"η�m�L�AaQC��U�_$dm�����L���=������tVB$��Վ��H�B@�w��㇌K�{׺�\���Q�4�lL�>+��C" ���.���(��\�ŵ\��|����s�J��'�y��	g�f	s��C�EJ֐&>p��~a`mruy�Z��]蕧AC�r|":�U�aV�q`{�xw�1���󧴨(�ݪ�r�3+ۖ��c�Ȍ�g �y�4?ƍ�%h�P?��1W떻Qcp�����L`�p�Q�ڟ�s�P�1t�|5ћ��eiw���|zG�K���yJ�L�Q����6�'��3薳���4��q���Q��N)	p���/��n�Of_� ������}K�M&Sy%F�ZEx�u����h,�#���~+T�F
^HC��=�H7@�A������0�U��#{_�(ᩢ��u�~��z�A�\��÷�F��m�������@�A&81K��k4���j@�M%�84�7uAjk�ƫ�op��Ks��V�|�Zg؎�&���y��������K6���r���)�&�
s�@��BUў��mW�$��<��_|Yt[��Q�!<z����I��U��
�^�VK<�&�
�It���N�����-�,��{�si���{8|&N��Ao�U=h@�3U�&����ﯬҷ6��|��)��F��ޯ�@@�@6�ܮ�?<}�EIIIQI	�榢6�K�J��흉�a�W����e��M̠�T=/L�O|y�$3�AD� ���Ax_���;�f��y�q����3�9�+%�X���MH7*C-UX�E>A�{@�V`����!�9��rr�obQ�2�ِW"'�pӥb�=�� �ȭ):�|��Fǥ7��ykQl��Oh�{3�&�����G���TbA*���H�Ǯ�@3��PU�d*��7�Ș���AD�+�?*a�[����>P���]��"l"aw[M�6<*� n��c-�4��+�h}�aPaI�H�z�(���k]���˝�����4�<�}���sw���X���u=����8a���zԨӗ�Y1~h@�����%*����<T��`4���$������Ma���R/�2y10}C�{ot=��q��x���aeu��8$��R�p��u��;�'߱E2���Ր�?���z_�>�8m ����L}��d�U$�ʖ�������<}��HٌXX��Hˏ,�h��f����͈O1��z�A���=8�� �����1TD
�a�����n�0�Eχ\���y�Ћl�)&Vu���M�̓�L��б�=@�26��	I]�P��E[�,��������dc%�X����K\@����J�(��n��X��.�4c!�2�&'gQ�C$ �...��_ڥ���!�}W��$|�~�v���U�A9�m�+���3�mV5���
8�Й`CA@����f�� �QSSc��Q!?����v��mjA�:c3Zb�kl����6��5�-xv��h��|�{��Gt�
�[d�z�]'`h�EԸ���H@WS�?H����;���c�y���߿�N��Ü�~��վ���_?�d�y�IUW#r����՝������S�(fO�Ҏ���C쏲��� �����Y͈{��MeSC�8���t��&~��3o�O���7).�ʫ��.��i�����2��o�����u5��Fg����8�A�+��fs2\�p���:b�sZ�ĉ+C�{x|.`l��'����'}f���QH�zG�E�r�&�%h 5P�,��q�4�=�/_Z��BzzD��^�SXYl�D	ߟ�����VR��m�b��k9�+����>�d������3�p����3���6����
�܄p���i��֍��˗���*�9:��<�VN�H��0d�&J�lX�؃[--!�[���V��p#gG`���#�?�],��qa�a>~�h�� �)3:��Q�`45�y�K�l>]����8��C}�O�b�T�g������xo��VEM�h�#֫Y[�8@1��ln�8��%��4s4�K­�e�w�eӀy3!���I��#y|�фUks:�����R
4-�jO��W��Om8 vn�.��2����yd��Ƒ�{���7��x�FR��+<R�+
�׭�&&7~}�η�>Q�4%��e��Z<b���- 2�gg$_~W���� E����/(�55�)�����{���G���MOQH�����::�9�&F��͠�c��<,����簋џF�S�+����,��);<���{5l�X�������Y�<�H=�^�6�H�}LyB�������Ѽ�A�(@w�~V��?��CG�M��HД�s�b8�b�S��	_G������b�E��m9�6,P,6�Vxlz&��7�O��?:vϰ3ǥZ�Pu)z�y e3v~BX��߮4P����_�6>j!�&�a���}h�xkS�i}l�GA�M�@k~$>�6&% is�+>�4�&����w L���}��<�0n^�w!0N�Q.&W}Gg6}����|ރ�;���H8W�D�݆!��0ȭ�k.zU&��ÜsVT��lK�n`��
F�+�:_4�Q�x��'�ƻU=nܤu����r�d�M���xǮ5ߥ�f��Pp�;@��C?��Y�QY��|W��ʇv<�،d ۝��)X�b3~i�B�}��|���˓j5���d�P�4
��&gWw\�@Uh9B����T��X�'�\�5�;o�&�х~}m�S#?D?v��)���U~��9�o���Ŕ�o����ڝ��D��v���!�JO5+���ɇ����_�ݤ�X�9��JCIa=��&W
*N�-l����� P8���7Z�M=\92�L�P��?����YY)H��2�����zVUTqb����sG1m�X�PT��n,{��c�BV�̒�ڟ i1a�����V*q}bf]�� ��0s�ǲ���?���L_��2}���j���G�-iu�/#74����c,.�y9ⷵ�G�f�TR�,�3:$���D��#Ϗ�������U�\LLP}�]a�3|(�E1�f ,:��(���6G#�����"*�x���K�1�p�oΌ��|���|@�0������PZƍ!ƍ�����V6����y24+���ޮE�Z����L���Y��f~h�x~1Fx�f���3/�d"�
���Ti�ӹi�>2����T��y�	��e�>)�y�A^�,N����~�q���](i��2���j��_��O2���vC���Jf��߮,Dvν�=���)�=<�V+�V�������ۯͩ|�}B��c8{9�oH��:�����h����\0%C�Y���ƣ�t��3�G[��eo@�i�_��a���t�􅘔��e���r��}a�cg� ������Ld����ʂ�1�K���?�D*�q��bb�|��������ib�h�/X�����Gl$)$����4�5�*=|m��^�a��T������9XV^\ZJ�����V�YA=����v2&�ym>���C��t*5�����b<�|!(D �!�q��E��\��êT���M+��ι>��+�]~��鵰����d �賣�v
���+�G�ر��A�"��r�y�h��~%8.����hh�w-���.
��ߛ)�Vjq��Vܲ�25B�oc�,7��&�N�<��B�/:��3��W��FA757!��
�:��Q󌘤B<�;�2;[fЩos��)�O	~�qJ+���È���
�{�5��ʧ��Cݴo����-�Ō��B�y~�:6\�̱-hO .	���3~x�m�0$\F)�ۓɹ�N�T��A΂[�̐2m֭��+»?4�滊��'D�����g[2����m�ժ��$1��nX�K(�\#􍊍E/�}~<�df/�4���&zxjY�3��(�8�Ͽ)���,�pa\u[ۅ���J��eP��5� ݑ��'9��/����c9���w�c�:^nu�ǵ,*�������HI��^0�jv�ea����R�l�sV���R�^Z9�yJ�����pZ��2??���Z��F�-����x���d�^�d���Y�B������g��d.��)#�����*��"
�x�٢]�݃��ﶎNp�Hj{���0�aotlLMa ƔLg�����������ՊHX���T�R�y~Z�����v��5��Hɟ/r9i:+-�\2��e�%NS����I��V�nLZ�n>F�F V,�>�C���REk��� ��ג�)Tp8��X��}3�ru����V%R��_>E���9��s��W��-+�yg�ݨ��r�z3	+FH�`
�^L�{���#CC2�մ4��n������J�9		'''��/�x���~Ya?���k�Y9�^W�FT3#�P�R��W>����:���+�T��J�4�U�᜕�SY�)�-�i����<��5022�c1Zd�T/�|�S�?(�(���a��<Z��{k��k�(y����g��ws:.=�}=2��
�m�umr���~.޶[i@1�}��+�����D$cH��f�I��Y� V;|t��T`�v|���)�Q``f�4X�v���Qr5�*�"�b}��U,�0��ֵy��)="�5��\/�!R���2�tN�����0v��/Di%8��>,�A8�f�	b���#�{�%�˗����������sPUm!7�[��iE���2򵋭�9�M�\���湹���1ǘ�f�E3�u�]��}O�~����4X�#��16������'��s~{+!'��b��_��?��D�Z�	`�C�>� }�;��6�{W�iq�C����UN$��/��u4̚��@d�k�]`V�C+Wc�k������Ӹj�&4��RX����V�	�^�p�LK����Ѡ㓂�2�azI�"g�g���e�U���v�󋋸��@��ύT��64>Q�B�3L�ʷ�4Ui�.j��|b�J?;�!ſ�v�(qRv#�D��\�=�^k�{��[T,Ϛ��O[�� �6Lw!~q�����+Z��:��Z�����S�qvvfv?7����&C'��+Ygy������H��9�p.xi1,��Ԕg���~�w��!W	���L�rs̚6�1�\��u9�n�'�kTd$R4� ��5���\>[ߺ�r�H�S#}�XO&��A;H���-77�L��{ށ.!���g���g�d�]\r�-�u���"�� �-���:����Y�\\�T<�J�z���6?�}ߢx��<�F;t��� ��;팏���p�rt��.��G��v]��A��R�&��-���HCI����֢'�O���ץ�(���C�������aɞ�NTٻ�m?>�q����s21�j�b<����L�_9%�41|��Rt��ml>�����-�go-V�r�hn���)-uM�c(v������啌��f�֥b�;�������E�E�^�m�U��o]�Z��ԫV����jTǓ�g4����(��,,���W���ϵ�;���=����O^ԓ�ߍ+��Ӓ��?�Y�*���Z�`�󭨤�;FG�gU��q�L�Pɢ���2�C�;U���ο;����rȟ��ie��U|������AH�L~+���ك��2��h%_;pJ�UM/�1<9�{�O�2����󉅔�9^|Q�܇��&����L
���b'�ǥ���?����C����d��$+޵�W�Y<m��۽Y�Ҵ��r.5@L�n<M�u5�0R��b3ۗ�t�g[R�1ë���e	���V�F��oTyC=�s1���FEE�;��U�[O�ȥ���l����x�����|��a���r��g<�"�{L5�H���D��*oCU�f�!�<KŞ��6F�]��R�������D�^����@�Hc���!�)������I�h7�}oj�q����	��R�^�L5KV14�y�YA��3቎�w3f�72�X�xa�h����������S��b�K��Zo�9�������0��͵��~�[pez��Y�Pث�A˸�ccc�Kl�KK_8���8���������c穋o+L��x��u�����)�(�)��;�t �(���ѱ:��Ҳl�r����}�f��4�U����0P��A��8��	�C����R�?�촫�4XZZ�Ɔ���m�R�0{X�O7�0��j��^(c�k�W��%WJIKٞ�Z�x��k5Z�.vCO
w��=ydV��RBBI��(Ԏ��re�Q����)[���}��H��w���}��}�3�;���c����qRA	u��m�5٨o.R:���Κ:���'�����;�9�Akp�䯖%����a���1$��"H����EC�f'�E��A@eAg���G�r%x��kP��V�K�"v]t���2_���U�LA�_���ƽ!(�u�,#�'���K˖�{��	W�B�'pߴә���g0�Y�IA+((�IH�����֚4��"��gg0&�J��H�����;�cQ�c��)����X8����W�|ۉ%WqI��\+B��2::�0�ĩ�cMW�
��k].</D� ���D:���B�L ���?cIk:]k��&����'ߢ8��ٹ����N�T�UC&p7]��}�R�͛���o�wXY���i%H!x]��wK-�� �n���K�6���h�Arw��z���G��=�T[�񔓓3,22��^��Ǜ#8�dzW] O˞��I\�<�W��كz�ynN6��A{�����J�����Zf���c��54l��e����Mn���Z5���M����i)S�7���&��r�9"�z>�l����u��NV*xy(�_FX	K����\n�	��f�ie^���$j?K[�Dv�03���wQ�b�|�O@��MLL���<���]S��	ɑ1����^��
�'3 �Z��3����a���ޡM���a�k��"�����Ty�+�}g���z1����n^�C�}?;K;�������
;��v4�����O�7�k�SSS�3�2'���xlf��?�K~\��Ā6�T�P�gb���9~p��H��Yt®��U�9��$��u��ݹS^��{4�!�Q<�e��FV����ߵ�t�DQʫ;5����2���u>������ٽw���{id��LLPw~�=�H�Yws[��� �tuT����C黔D�ҝ��fjjqj�D��t>Ƴ�j�F;�һ'�3rTox	����T�ۚz'V6��,?E��ή��0��-FF�&�;F[��EE�Lr..`�Iڝv�E��fJJ���ӭ��~֢�'������z�Z�`%����K�OVS]��xT� �;�՞YU�i��+��y1�����'W�tOS ��+*�\~Z�14���F�}�|R�f�U�5�I ��Aͯ�n��o�`�uss+���� ���F�>�G@�N�H}Ѱ��,�*�-ɍ��U�{*hI�KӠ��m/b�R�d�8����?�O����PU�y��'�'`2����]�������|6N����쯤�ᥦ�[j8�t����$�BG��]���]�ʥ�������K����@Zk>1�#�+��|K��^MM�x�`�
H��-���
V�z'-M��w�ȯ��m��)��4GF���?{�?>z&Bt�H�A��ѓg�W��;��}�߯ʸ�q�綦�VP��r5��^"q?�f65�a`����42�6�`ў�D�B�p�x&��	�V�ql>??���u# Z)H��H��YA�oy��F}�@ɹW���$����c�����z2y���j&��1��E)��z��g46�v�?��<��@"E�xnpIs�b5V��o�ߟ�q�q�?7�����։�e5+V�g�Z�S�̷c_c=���!a���#�������
�	��������o
\�!C_��Q�pڦ�Z�����G�0�e�@bS>fhb�߀����$|xx_T����p���������(ơ@@BBj6�h�E��g7��e���_��'-{DB��<I4�N_b			�rr x����5Ϯ��-G:���^`��]'u�a����	�����i>�(�F)J��e���@s�������L��0`����n�������$��\x`���p�qd�m(µޅ�M~����#�^��tZ�Z�:�
�ؒ�j9C4WG��,Ԍ ~ԫ��0�����7~��j���)�4jhi���z��M�L&��xyH�---aaa]��e���@B��QR�uW�'�h>?�-.�����2Ɂ� ��h��_��+ՐiG��366��%��<�����+�
�y�`#�x���XN��RV&����?�M�O�a`b��Qy����x�M�O�(�Oa5���˙�x�+��z�$�`ih�SoL�e׵���¨���3��x*5�ag���8�CB�H�����G&�F��A٨�d�و�X�I�d����3��*XAvj٫ ���r��&u^�͝��d�zF�?�-����"#k���<'����#��k+.FI�[m�����2�F���H� (�	V��GS9�ZZ>��S��-E"�c������|�LNC+/?Mڐ�����SW���>� ���Uȟ@,��Nji|ްzp�Q�MO��o7<kM�d����1R0��{���ݾ�33������Q������W$a8���k�9qr��v<e��DNn��A~c ��w�LO�^����)����5���r�n�v����ݫ��hn%����n�+J�v����\����Z�ձV!��`�ggU��ݥfg2�!B�W��oT~SZ��Pu�on1'$�qp'un.��'қjM���q��{7K;��w/@��տ��� }<��6���!��鱣:]�����	�EΞ��A�n�6cQ�̂3JiNKl��w ��f�@;����VWA'���뺇�������"ï!���K�}�//ĴFќ��2���%3@ �{i��&=AM����D�iY�C�������-5�dfg�����E[����#�>��T{?8��{>߳H|'N#89��OW#̬����$�и�Ug�WWG�}��Ł.�Dd���"Co;�55��y�l`���r�5J���٭�^\f6�o*N�Z��V%���ކH��5�����x�a��g����+�	5l��bӼo�!���rrS�����Ҍ�}ir=! &K@d��Z=dq`�t�'�37	��IŨ��S�5�	�7*�@����P���'UK��ӂ�j`��?�+52?'SQ��4�؄]�x<Roa�/���h����)N��_D1�g}���؈�C�:��Q�pO�[���^�2��K:}�o�-+7}�ԯ5�޷gK�*Lb%�6$��^@@�u���� [��m���T�(�u���ա<1_K�n�5��%�S���M�{Z������˫+ЦP���H��g1���}�;F6�J.to;���Az^e��X@�h�}�3M�;]�,�Ή277�����rC�w�-5_�c>�����1���\b�7�F�g*O�{���M�� �'�Ղf��/u	��s*��MP��=�~���*���d������1}N�M�����:��u4���	"��UX�X���@(F��0��F�� �A��p^����)�����YPe�BH0�����aXF%x. �W6*��W�ߛ�@41�$�䜩�tJ��θ�R!E�j池#��V�����+�PT�o111}�>(����a�6mGb���g��X�<��/���8q���o����)�����~�~&��`�w}8�DNN^U[o9vy�L̃�H�e���B���1�?;#V��G���b�� �?�p�yq#�A[=0�GG#�o7Gx���Y�~��'�,/��V>N�m>��a�KHn];�iy���z��F����O�.펦b.����mg�h=���X����0��������r�ި�@#sʕ1� �\cL�m����U���N p�g��� ͋9;��^�-eXf����(rw��S��{���p�L��pU���輢&ݹ��),&��kK���;ss�9�v#���5;2�>����E_�&j_	�s&��@������
�5�����ѣ,^7�����+j�s�"p�'d'J���NB��G)�=O��T[���C���r���]����w���V����lT_�+???44����+�JiI	��f����.��xA�$����'�F�h�d��?��,���f��]BB� V����6Yh�N�������cT�#��q�=�e̧k F	���EL�o@�XyU��H�C���?وV!Kl0�x��ܦ$''�b����̌B@�&�F$}��l�����������~�ʞ��b�EB������>!��q,2!'2 ;	�CZ���a���T3Cz�)t�������Q(U�nT�.�_���j.�~���`���Ykuc����Z�)�������0.E55ꩶ�ҫM�a�5�M-��1+�^��}�ǈm�M�Řw���x�5_�HŔ�6컾������|�������W�$ �?T #3s*_7��c���'s�*�Z!�US��|�Ӑ���C��>{&�bK����>�����C�$k|ZD��5�ԅ�����ы����7rUп�������Zz��uzz��T@43���C�ʊ�B�=�K<M@o\y�T�8�h�~[W�F%U%fxl���[6�aW���n/g�5k"�;7��IN�����54��R��a�W�J �p�Y^�}�/��u�?�=&W��(yw�f=�#
'��
�F�'dfV�w�9��D�aj�r�z'i���#�
�B�Yg�z���97�w��v3<2r�M>\��CH)(ƒ��/���X �5�[�XC��D3�Ӌ�l���(���U��xy	100R���!���FYX��	�����M��1�]W���T0�U�l��4��>�^̰p�>�FD��J;����leq~5!h���yV��	Pr��m-M Ho�@8��������fY(��īm*ۼ��g���t4���� Ǻ �ul	*�-]�[��(��@��5���JҞ�^�yu�; �|�fe1j�	ø���>�i��gxc�Z䏷*@��C�@����i9���~I@�L{4�T���~CB?��K}�����˕�V����-��Xɪ��+�;�T�X�]]:6��ļ�rB��h��g
'd	�O�~!������H����6��C}]P,F=�}�2��=o^Tt��*	�F�&�PP���d�L]�pL����ּ#J膖_�L��:�H������蓁��"�@w쟢��uQNn��)���t�_����0��V�����?��,T mjj�M480 ���QUS#"+���BO��~M�����2��p�,)��0��g��G{Sq	T.�nW�RޟG>Uu������n��I�\��:V��5����F�8%�м���F')�F��x�s�2���i���w��TO�|�nڏ�4�Վ;�����> ѹ�|����LEEtF��?�cYlc�}��\ɪyv��5��cJf���_�O�P�||@�ۈG�;��C�>6 �HN�I��_]h@���5�1ww�_8t�2o�/�&��0�#��A������o�flfb�� s�;�")/�:�(C2�-�k
Rt���]��UW����Tf��O ��N �ˤ/EL�ԉ�u&�t�!kjU='T�8\����� c��`�&|����\�,KFF:V�߳R�L����� ����*<�w�������J	��PF��?���,�.�c%h��2#���e f	�jB馕�Q >�Y����ٺ��Z��U�6��ᄍ�J��(Nl�)xփGRS��|��< 2�e�K�� ���
>yrB� �ɿ��V�����0w������8T"n��*��UU��tB���SM@�6ק�!�>+���޼���..����)��Ԧ��~���]���knݿK��!""��fo>�9N���f��[�ds�?��u'Q�^>Yc*��������gQy������L\ZZ�B�%99$�|b���%3~1C_�z����.VTT$dd��3�`Kc �ltd��x�7|�;��	v}a��~�������,���=�YY��dD��q��T�q}��w\&>\LH�
�n�' E��/�RY�[gg11ʣ���	��&m�=ic�Χ���D<������Ō�����K6�;�o߾U٭�`aa������mɵ�l�+�����e_�8ǜ�2�g�}� �t:�}H^^��e��M�l귌���a���f����R����~/.�檝j��[����/OwO�#z�W�R8m	 -����&�B���������KMME�&�OЗ� 
�'p�7���
T&��>� ��mv����������L6�����V^�y��������GlFFԯ_T}���rFGs�'����p��7HG��*��gD���$c^7��e�����'!�/�rC��+6�����m����\ӑ$�{Yx�N�bݿ|�r9A@@�A������9G2Y}�X<��c���V��U�{��K[i�-9���QO��/��VV�����THִ�:���q�/��$��A��������1��[@��Y΀���Yk�D�������3E�Φ�}8c�vW{;�n�M�W�� ��&����0�~�#v�b2`8S �?�����I{��N�\[�w�v)q���]�6� �Tn"��?V��ߘ:�߁o�OL�fN��iq=� 8i�=K��/w#7�9TDDDU6K��ق����,�4������&��+ ~Ӫ��..=��h���[��߱~/o�L� �,v�	�{�'p�I�vVg���S��3�՟��&1w
&�}�������Z$�9��+]���^���Z��o�YY����  ��xc����krI�V�O�#޼��@*�,�=��k�I�&������竉���J�O�txy�l�Z�,c)u�#DDE���eX�����x�OI����i�Ց����1����r=�>�A��9G�NS+�F�xn�2�GR��ŵ��W܏� ��}��r��"�����?����<{�b�,��H�@�# ���M�q?b*j���(|�*�
X��������z�jЖH�V-,`�薆jcc(��� Z��pi
�������v:��}�jzp������biiz�L鼢����T6��#|�n?��u���c`�4���X�\^��ed�J2@�m�U���S�$��%�ĳ"��q%��@힘�o����N���T�oz3�i��o�9�G����Gӕ�wg�*Ys�a``��]��++G�k��{�����1 ��@��%'�j������.RA���k�,�!yՁ�۩mn<�#ń�>O�]�e��I��j�����M|��Π�\���LaL�����#�,��D͂�`ۃ�����l ���������b5"�����������m-mmc�@����cb���9j�{���H!�
����A�MODj��:�����Ś��M>�/�dPp�1�=Z@����5�ΛrVqRAף�@VڙN5�N��	�h���-!G��W�1�K�F(�脖q��g&E�YX��2&.�o����c|0��"�'���"91��`:����)V�!A�~�tֹ8!<*��&���L�^+�Z��$�mW8�G?��2#% �����=��%��Wa�7C5K���MF B��ͯ��w>Ȉ�%M���֯{X��O'�����Y #����[�D8 [ΕV[/0~_u� ��(=��m;���b�COW;���۽�����A f����ǯ� t���\\�{v�pp"��6��L�v��T�TV��?��]��"]�t�(]�
(��HH���Hww7H(���������}߳�]뺀�3��'�왇��K-��#�>N�ܐy#J�����)���H�Mq���x��� �f0(���%����J/R�ӛ0Q<b��J�Y,J�w��0���گ2�������_f-ƳH�55{z�[w�z�����O�;m#I��Q5%?R���z��ds�l�7q�]΢d�Nv�����Y���_�~uu��cC���KD�0��_Kc���C5�Ƌh��.;��������@�߿����H �V�?��� �z��������~�p����*����-R5��:�8�g9yybo��z{�	�8�3^%>?8=���簺w}�HYY
@���������c�Z_]�����A�͍//??5;���(!!!E"{c��Y��t� �n�+�\�Sl>�v�ݞ�T,�N�@.�|�133;�q�����J�]%rWKEI�{��n�'���+��ǙKh�����կT�Ҋ�7o�?���-�������������]�\�LH5Iw���eX�N����w�qq�		��g����c*�\�:�K�'-����>A�[�N��������t~�Ԓ�Xq<)���l,���YM+ �.��xH�I�@FQ��eK���ݺ'�TNAA�O�|�XQ7d	�FD�}�s�81{�F�%=>���Htbb���������}Y��ŧi~�2������Z��?(FR�]�C=��6��*�uߙ���f��	��?}}a�FLLL�$$�@Ez�h-O���%y<���ZZ\T��y�]�����i�Yz�d���ެ{���	�yݎVQ$@  �Ԟ"�-�9n.���+|G���"��"��s=�ڗ�r��뭹9: L0��rn���Q 	�t���N�Ɔ)&	,77�(Cu���}Z����Q>?R���*��� [H�HK�Μ.�~Z�S���uNACK�^��'����(Y:q9�̟U��3U���G�:��MOk3Z�6y>� bQ�x��v	���1��?~���K��7x��������j�y��	����\��O��#Ƭ������P�� �J����� ͋��A����l�fpd$��
�ĵ`ҥ�&�L��E����K��Bv>��fq蚷�nP�Z�"����V�p
���Z��������^����@Wx���:n �3��LLNj�iRyT���oim-��4���yyCoL'KW�K���H���}S*'�@@��f�~'�NN�I���&\_NN��@���:������X���R+mh랚z8??�����l'������H:r�f�}gK.r�!���.��f�--���#�9H }�8�L~((`�������ȓmnn���Q�Z�0#s���ɦ*T�7S�|b�(�����p ��AZD#�;.L/����۲�@Ů� jgǩ��
$$�45����T�|�Aի_h��LU����=����0�V+?#8��?3UW���Y�###�3�ϒ�g>� ���D�`me��A$gd����Zj�/B��"Im%�|�J��[����[1.	�Dؓ�AN�������># 2�K����i}k+��s��֦�6���CO���z.��մRiR���J�͍���e+P�KKK/t�z�S�&=x��ʠ�j��@���=���������&���'������5��=#�C�(@�9�X��ɠ��}���d�ϟȔ����eeQy��(�_�����8n���ֶ�Β[[[k�92>��_����"!�|[k���Y��skl�0�[���*�%6��R[�~�Sl`�3z�\=x�k�����b
��1����I��&�j����΋�H���\��H�8|g,�����64�mONM-=�r�=����H5���*�� ��L��ox�C%ܱ=Q\�u�|�;�����s�'x����̬:�/)�ԚĽ����ȯ��z��A$)�9N�ѝ000Z��s��0���u1�%�o�w�]��k¡edD+6h���u��������Yd�����|]���䖫�]'�����T�J�"kjj8͚߿���O�$�уSn���bV�QF�,˩2)K*W��)����(Ł����[7�!�q̚®�V3U��|�F�}}��x���{z�+ 	�'^=���|[zZ���@����U�X 0kJW�k?~����YdxdjEDBz�ԗ�2��^ү�ϭ�%%:ٞn��7���yuh`�`�DtBB��i�s
垤a�BR@a�q  ���	z��Q��u,���<���Hţ��
@���+*�6k�%edP@�ٺ�ȀO�U}�L���v�ʡ��ࣛ�v��߿-ONC��;�<�A$�y��k�}l$���}ߐm*H��Vfl���i�It��S�jpޟ�6�1n�#�{�ϹԀ�F)>ߝ!�d�9Ǘ�x��	x�w��I����K�7���N�b���� �tU��������$@�q�g����h�����O����ё��@mݯ��@��޷��P��j�B�9���D��u�/� �z�}a���ϟ	*7�l޽TH�p �`P��wP���6j��'{n�s��U�#5���^ ?�h��.�mO6�!����YĴ�R!�HNݝ�?|�P��qmmRUՅ{ff))��1�=�_�|)�������eiy��Χ�bBaM�+"<��ͱ��t�fl�nnnr��� B��(�����auE�o��o1W!��>Q�\w6�����q}_����/�uEMC�����jq���p�^@�t Y���[������n�ק&4��u�4-Ù�6���i����i�e��a��B}j���H�is��Dt���u����[�<�ZVY�Yc��a=[s�ӵfxs鐑�u�����G??xBBƌKccD S ��x���Yu�����#�y�@s@�ݕ<��8n�$�Ml]��|#�;S�P�B�و��K^>���W@W��������bbfn]9��EU���~�x��."$M��(<<|�x*��S.�m�.TuNZJE%&o���!eF#�!gww����hӂ�8B^r�ݢ�r�P�o��+��h2��֏����D�}�	�	soZ�ڗR�A|rpq]MT��bZ=<_^^v/�=�.����Uj؉R\m5C���_ށ�DU٤Xe���!2�F���%1��C����I�NP���iK-�µw�v�P����y���\5u���ii��	͗�^�s-Lh�[�z��$l����WY���Lr�N{�p���k��(H�)�K��yl��$LNNN���m�DK�?
 alc�|~�ač�;#�o��f͔�2��3p�7���:~��(|]��ݾv��b(���r=2<\M6r����VV_"O��@��ǬW��H.���|��E5�u�~��`�phye����Kh��祮���"O���tg�l�9�`ӭU��L]�,�((���������rg������������,���l	�z�k&h��U��|Q�z�I��++�%���u�M���gM�OEE�{@�L�]@�Nx���h�Z<����h��A�|��d�rtL9I�[G�L19;��ɮ)s;1��13���Y]��8p'��8���w�s�Y�^�i��#pٓ��l��O�2��'�u03	�^�;;;����'M������5킩Ǻ>�M7�ކ�����>۹F����	�/��;È�j�{�]� :Yy�@�i����v�y^��=U.�G������@ٺW���
�Z�_[��+	u����A&BB�spˡt��L������'���ަ����t:�q��z����R��iB��(����lUp��R��ӟ��u` ��f^�{��^F���(M�<ۙ�=kxhe���ρ��u�4�,�� m݋qH8R����t8~�����
��*�C(��'� '/ �����珧�� 2�Ƴ��/��Nx��}��'`F |l���( <WZ> R5Z�B}�饦C4���¦H��|�7���	�P�����3C�-��B�g|"��ıߩgBL�Q<AD�#I�$x݈�'��a�I/i����d6���
@ޮ�e��XF_��b��6h��V	]��y#4�POm�D������Z��X�`888�B� :L��2�FT�������aa�|��#���H{�^{�S��6v�7�����ʟ��X�a7D��_#���	8����3э}��a8��~N6E�ÿ��)bma%��~)!�L X���=���_����i��»�e�VQT44<�ɼ�oJ�&뜘�_};i�~���d�;yZ�L����.0�@/��x�A�F�(�F��/��hYB�O�|G|��j>���דM^U6�����B-xM^�7��2���@��7E��~i�{����C`�KJ8�`���X����$���).��)d��F��()#�outt������p��[ckS�v%
�=��У6���~��A���o1���rBb�����B��H2.cT�i	���">���I ���+�Q�A�����r�b*����'Pk���~���F�w0nڞ��6��&��1eΖ�q�?J��|�zvVV���;�lA>�!c�A)�X7�1U��_�kh�y�����l�a�	S=*��� &&��a]�D�����թ���-5559�R_/=;:;��+ �F_dЬp��-����G�J���������)R��N ��	sr���6?˵X��+HЃ�3��<���dv7�ҿ�:g�Z�����|����f�:3��4�QϦ!LU
0�NK��wrzEͯxv�k�t�(�W��ApȢ�>t��e{� ���&Pٙ�g�VʭI9�?��6�����4lqy��ؖ��h.�v���3b>u&&q]]� w�8	SVV�Z艩�'a�LXsT[by���|XK)���WR��;�uq�^��*�B���!�+����duu�.{�b���`�� �
h�¿�������π__T�z��8B�"�-��:X���r����D��@��F�n0����i��4x��a<���-��,ǡt{J�u��y{�KH����/�zD�<�����0!11�w�g������1xU�T���"H�<���~������G �@�zܻ�c�U�NN�aa@`.ܗVW��v�h_�=0 ����W����K����Ah�W6Шb,ݖ�x�u����I���}I���	/�cie)qT3I�����}�%����������iii���)����� O=�&('0��*y����6�s��y�����I]\�`e&ߦ3��.,�x����7x�.$�FFF�[���RPP@0O�O� 5'@���}Aa�����4����x4l�aO,���$���13�,����� ��������������J�ɡA�@M- h>��<�]ң��!������U��㞻�a�[=S����'#������vd &r{��Zhג����B�-�4h%X����|&��ig���������
����-�������l�5�B�8���Xn����ǔ�%\t��Q�{~��|��(^a׹�A\�?���UV>{��e
p��A0(�4�?���\z��9..����������i���/$��Q�W��U^���	�l^(�z�0Q6��B;����	-�(	��H��+�9�y����D:۝)�-m�v}k�i����E ���á�������H���O�x?�xԥ0�[��2W_���D������P��e�ꕺ:a^^ާ���-5�!���ODQ}��XY�7�	U���q ��g`�Z��B����I�? ���nf���68��m�"�	�e���tt��9	�\�%bqri���ed���b�ճ�D^��+���[]���'<����?�ɻ�Y�`m|r2��΄+*J ?,�G�y˴X�����Ĵ�H����,�'i�}=	B���D��c�^_�~z��۸��i���۟�ڵ���1���h��$���~*��Elu(z}u]�<��MH�"���Q��D��z����38$��6JPeE<��t8M�X?���{z��+��m?ݞ�~���Z ���������,��L��zz������E�8�o�hU�[�þ�(k�o�iZ��1<�Q�����N�_�76��K�mT�� ��(������Ǡ���h����9H07��y9L��uRb����t-��G���v+O:�*Z�_���@�s���#����iD��<����dsENN�^J=�Pj$����C��Z�kwr;�e^hD���ޯ}4s�̹��-E.HN�����-φ�Ѭe1��!����+7��� ���{s��g36�����V3@��ݴQ)�Lc/�;n�	y�� ������^�����;�������ӭ1�7��+[�Q`�WZQ�$_��J�L�G@`�\x9�����di���γw��W4i[���*�v7���i^�Dqon�$&]6
�n�a���I�ku����R�['>�ҫs�j���'�����I��A�Q�g�3yEE��/1͘�& �\���W∫@��s*�kv���gܭ�1��2�8a�9-��`{���[pZp{W�
��F�$�[x�ِ`p�jIK#�D��ҧz�^m�T��뇷���P�;2���*}1�����9�c�'�]�|�aa����oJ��s����C҂Q��fʛ��N���V�(�~�
q����y�P8�a��O3.^���h)҈���F�1d��cѮ���~�7���p���}y���́Ć�� �k?�����Ӄ�T��h���s�H�.֫�Rz@s�����ά�Ob#AX�|8~v��o�������ւ��wFhMW���eB�$xxS2��!å^��f����R�����a�`
�U:e��D����e'��RR�3MZ�#?��N���}�t��"�	�E�6F��eZÔ��������� �u{-K�ʃY���wSddf��ͅ�/��Q�Sa]�̆%>b���ضmA���~�-w���P	�I���3"�˞����vLl,�K	�����m=O�x�����X'df4��J����$��9��*���?�3cT[��rn"�?��剧�
	^m�#��ni���z���~��0 ��e����ܴ��[r�o��b����뼷]^�F�a#�>��e�V�:e��5)8�a����|��V���m��,�b�w����PzP�[��B����B����4G���h��1v©[RB��(TB�X/^D ����Oy�ï5������u�&�+L��T������(V��7M^6��t�� �]�����E]pb�j���$�����JR[��z�!$I��p�g����kDd���F�c[c�ˇ��T��T���lOȕ���G<�� ^q?�Z���e��1�9O��.���׎&?����z!/ϪOn:]������8׺�٤��9���V+����r��?�\�K���jl�}�㦡�x��;#h�ڦ�?Y$��SC ��#<s5�)����C׫m�jD�.V�jl}���m Z;���B�y�m֝�zb�k�"�D�V���P^��kY�k�k}�fFs����4��DB�}���fo/D$$����V�������$���rZ���/��@�y�G:T����jzt����6��p)�vEI��Ͻ��h�5f'%�f�7:Jḭ�1��vH2@�D��-�wيɑ��Za���g�G��g�_'"�K�H�tޣ��~|şK�2ɚ?	j!��G0�"�b�]���Zt˿ޟ��Ķ^�����l�+J�x�7����9Y�R�\�V,5��LL��g���+�{��^u7߅��D.��K$�z��lon{%�'��Jz��5�zU�K���U-���	b�疢`�(�ʫ0�s��	;�Y���puTB;�Z�֊�͝��������]��B٢�(�Ω�I��J� �)w�p6�#R_����y�0Db��H.ě����,آ2=)�*L � $�=\$ed����7�31�n�f�U�Z�J��I��_���\�'k
 Rۙ*�΋�8u�Jj��00�?#)���W�O�"O.����a�B� <�9hMqy�0�Z�|n5��k|!Hq��BdP��_C���,�Z�;��HH�����i���)7�b:f�,R����zD�z'W��+KATEe��O��j?����&����a'1�q�'�cӟ���U�>TTT��@D��^�sY�i~,T���q�/R���N?�)K��5����XQ,rq�}�%�Z:w���>|�1�,��oII	�̩������O~�-j�ޣQ����PV�m&��ߞ�ں#㱆����H�qi�� C����7ӌ�rG�t�?��x( Dh�S���kQ��?���J�.9��;D�q�]Kz�ZZD{Dd��#��n-�@����e���ɂn��XA�T�ٌ�(���[,�j���K��K�3f^���oཀྵ<��/�[�֥��A�ʮ���za��]؜��z�>P\���KT��/�|�ZZZ+vi�36ͅUs��T��˔��f}������NQ���*o����c]����(*���3׻��½�J�x��n��`<ו��=(��Nّ�*����\��X��QU��}�=o������V�4�?�4��vER����o��lI)�m�X9��ͥ��~,d�ǭ���4�!CC� Whϊx߸Bu�����{�O�{�m�n��		������ѣGP+���}�f��U��-e�Z������=@#���7���]o��ٶ'f���r?�)�ڟo�q?�k���ʢac� R09���T���P�E���pC����'4��K�|O-�_U�6�b��HJ�@�S<��*�|�B�*Ѧ)dxXE��z��?���9;C�nG}�A�g��]��̊x�YhW�f"�jok�$��.�a��o�i�B�U�����ק][�ͮ�oZ�b�N���g.���T�w�8� *�F� lu��!��r��~��$�^�ZmK @3Ue� l9[3����8���\�s?x,��n<n���-N���I���^n�
��"����^�:q�j��o��s�U�~�(��z6G�{�$O���=}�? x���j��Q��oO!O�ں��YyY�p-���۳;;�AW\�__�[�;����E�p�bШ)h3J��%�=�.CU)��k����n|�p�E������B�ӹ=���2��U�a�U$��Py�t��M|�+mT룢�n8ԦϦg_�D�
l~uM�]��h1ٞ����j���{ͩ�����`�#6�MR����&�*$�/�|@�Щ�b�r��s)�Y�6+T��w�@@�,q��mK���=ן�_���,�A]ŭ~H����L Jހ��zRƌ��D�ٙ���ʴ��Ď[�hP�� ����2�.&.�/%r�^��^Fp�V`�ɉc�L�cQ�0KO_�S��1���s#���g����D�@bͬ�y8:r�����}sǚy�w�%��R��?9�$W���^)�tN���]��T�G�dg�f)8�gy�d\t��Y�#�μ���l'��p��U0��IH �v� �s���;�����Գ�ru�پ=�
c��?�
����f�3��������#�� ~D띿,�f+$�B�P �,��"����zQ�fk��[���9��/��<��Q1H�4�.t?_ �QPh98p���NCi��7Wט�B>m˰uNniiLf�V墊��7�h��+�ؑ�b|�UX7��Ej��\����܈?
���'ˉH�X~�k�Y>���GO�
�\)[�b����n�K��e__��d:�DO�LJZzy3;�爢��;�ׯ�������2ӂ�>������������ ��%#{��|i0U��i��mU[�q�̓#�`w@���u>���̌�.sҦd��B)���`bOhmB�@�/��4���d�Q���7�"|�c͓����R~��^�*�|�(J�w&�z����g��������\�k�HJV�5�i>� `	�Be�Ȧ9�c��J�	�E����|.{��)B)���\�$�@���݌�-(`j�����E�c�[y�0����}:�h���.O�cE�l�*��003Kxz
���LGCs��{͌��%0�s?2q��5�Cvl)[��ث|��P�>3$�����~{��az�#٬�3�� �����x"����8��?�Ĩ�}�仱a
����lMCK+�\̳R�dј9��8�l����N�g�o�..�(iyS��s�̀����z��L[]5�d�s5J '�f��s�t��kiS��U���u������CM�6�h>��H����
�����-���;@$E<��
���ט
��8h:�"CƑ��M��V��9����"��D�.����1��-�_{�p>�1�|0���}� �t~���|Mv輫F@�ez�C�!O~�D��$�Ԍ���Pv��k1Q�Pm���I������>�x�k�����h�_X�f���n������J���6�����ꇇ�9,'9�s2Q�Nu�S�P# ���5������n̥��u�[�7���<>�`��6{ T��q�ç�Sl���a
k��g����R�ӥ/�*%|)%)9�W�+�9[����+DQg����������<�!z���Qq�sͦ����bU��7�G��͆�<��P@!��+�Ais��99P�&0�b���*+`����A�N�z����\��G�4�W�OnNF�6@�(�J7D�0����8�WV�@�?��fd�+{	��
2C���3������Ctl�? {hK�A1�o�
u�ixx&���Β��+HgသmL�[�yi��K|U�g�+�(3`�L�� �f�tD� ��+K�.3W��
����Ḩ��q(�a3z� �j��؝G���� з�P��缽	��+.
�Z�BE7���Y\4I����}߷G�,~n��bbJ*(`}�����!il���p�d�	�����N���1�y��覌�lh�UVVV�,7=n:P:��K�*�z����֍��t�.i����N�Xe$�����A��=�4��E6T�������9I�7"����[���q��:.�o�>@lllLMK+�K�-��(��^7�i^H�>��S����ik2@[�=6�{;��6ҙ0r_&p�����K�Lqy^��F����;tF�x&�v� >���t���B�pZ�[x��k=W��L�>��?(8�=�ٿ��u=�� (��&�)����e�T���&K�JA~�7�̙=�?�^R�����x�d/���d��4wy�-�+��N�0��h4Q��7P�R2���2�lP�X�8�aP}+�U�G�����S=~d��e�+�oͩ���R� �߂x3Kx*tS������a.�+�e5V��GA��\��}�Aw��~���tpTt�t&R%-_��6��퀼�`���XU�/����kp���=$p蛠Pw!�������G����ƌ����7������:Ӣ�ArI��w��UgI"�_�|U����s�k��;�7.�?f8�&5YcG�︑�L.�=�^_�N���T#Ҙ$����~�3mF#� }���.�Srr��bpEL��Cת������SOe��>���1M�5n��oJ0/�F�s�1/�">��R�3�kǍA�z�]q0x�qq���44R7G���5�{�d������ �W��6��S|뙖���̘�9�����O��a۫��m��Hi�3��@g�:�u�����b�K&*��c�����¯/�8 �MJ����`T�z3U��@�&n3�6] ڢn��}�d����A�&�Lڅ��N2�['�Zl�?�e.Ρ� <^ٶ��I��*�� )�1�?�'+��q��U��N����ݮ��������(�d2�F���f������tf�v����ŗ~���M~���wx�'���������ӂ�)���n��^�A�R�1hNKKK�����\��}I���쌌7;���U �/}B*�Lk��x���6��7;~5�͗6/���|��`5�u�v�ä����.��#v�+t:���>70c�������_]]2CōS�Ό6���3�Ű����f__X%�p�s��kH._��A�D0�X>ÚH-Ы_s�vd���W�7}Ti5C�C�9	���p���z�>�t��V��{}����7N��o��x���5�m�c_($f�+���zVI������	��y�]�X𿕴Pv+�vI���@'vL�����@?`\��V���G׫	 ��jؓ/)H����E�丟n�R|�ŃZ����]T>����yx����������/Gu�r(:�jb�7(g�)��{�����(ŧB����8��h��� n��320@���L�x�BIC����{#%����R�5��|.�u���c��0h���F2g���8}����k`�+�Z��\�5�o��[�@G��*'p�- �������X��-�|h5�#`�I�t໺���b��n?���[&���ؓ�$��**��@(M��L�3"M��LU_ѹH�BP$� ӧ�=hS��9ΘkLAvCj44���
7����9���)ejtR��s�2�9Q["F_�D����˜*71����ߜ+��lXi����_�6��O5MČP��Ms�>��#BD�Zڷ�T@�sݿ/?���4Rk�!���x�ʊ�(x���X\|S�ҽk��c�@���ZzVD�A�H��	k}>�ܹ�v/�<��� ���"�3AEjh{N:H<^���ie:u%%ߞ�'F =�e�֑�uD
f���Ӈ���g��N�E*��fC���p
:��v�o�Kz��Ba|�������H��Uu�L�h�P�2�ki�-n�tg�b��,b�q#�]%ݦ�P�;ԛ�(��>$d�ӎZi4��M��|������L��C�w��I*��_+��g���Hx��׃;3sOD/�!�{`@S�x�����˨5�[���7Φϊ���~V���(s���/����W0�w���4��ٟS����\�y=>~�KK��xp|ن,��7J��EY�����P���S�����϶+��<yթ�ޗ5N̄HHG�D<�����!m:�%��Ct�Wf������*R�B�(.�p�,�D�!	�?
UP����bS�mޥ���n��<d�$%���YZ�~�$E�E��K����^��C���KF-��K!���Ln	��ny[l��]h����]tp
��j���`��jSD�D*���������Be�2U����A+cI�I;�;�W�!�|���Ȕ����E/7T}��' ��F'�߈�kko�Va��	 H /T2PM�2�8o�'��������d�[����XZplA�J�C�!���Vj���^(��}��>9y8�f5Æ��#?"2r^B��2D9�"7��>miRa��\�R�o`��0+e�7.�0b9r	Y����y�I���%���|��]��w�>� SA��Ӥ��Q0}Q�L�,�HZ$\(��9�h��
K^����<�h�0��K�� ��CLRn�]�մ��%��4Qt�K�{˩a�c���"�XB�	�0	�P�NԱd ��O��K�����D8f��	*���W��+,B:r��>}d�-	�33�?`�:�i�$�i����-G �^���Nl����}�nZ�����u����	�]��@׉ ��o&9��y���"	#I�E��Mu�4�ĻG,ǥ�a#��1"�D�|ȅ�H��4G~��*���n���{���+��K�y��ȋ��i���H�����^�$�F��M��T��g������ �U��6ud}&�w��a&0D��P���>C2�`[du�b-��`ڢ�v���a�@�%z�7u$O�X���;�85=ee��=�ڋW������Dl�{��t��p�-:i�"h�g�Ch{�x��J|�
���s��n���/�ŗi�f�AEZ���hJ}���B^���*�g�2	Wރ~���;D�Y��H�Y0�8�E��CC��<}^GW
t6F�.�.�uy���Z���.�܊
50�RP߾݊�:��u7����sU��S�������I�5�p��آ�T���K���=�.�'�"l��	m �
�9mh�����������ve�*�>I"��pb�{�Z	������.���-��:����;�\��?�څ0��b�l��l�q�(�
M"�7��p�Ոpl�j���-�.�B{�.܊��0l�I�78�ܛ41�N��4�<��ňe�|ˏu^�����'7C7�n���ΆgE�A��[=����{
 ��3��#H[�{��H���2�5��˔{ܵ�i�yl�*Qeb��x�0��ΌĄ�+"cU�?3|k�����q[�����Ayn�H�5�>��J(�܁*f[�T�����2{P���α�8^�����x1����1�$�wЅ��'�Ν�w�nFl6r�*7M9�2�\���g����K�+��,��hhh ]�HO���D��̟DK*�d$����[I���S� ���=��#�����K���TmX�.�9�L�K��M51���b~6x`'j+�x�3��t��ި�E�|ssc>���,-l����=OL��z_�h�g����A@	B�s�p� �B>��\�F�V�s��Vy��*a%�x��s_�WYj�`����K�QD��i�?}��U$�q�����,f�[�P��y�����,h��/�=S@�X-̸B3�ĝ��2��}��竗,��	��_���u����6��/^b��ֶY>�֯�#{fP紝7.��9:e���ޣ��"�/uB�ؕ�_�8���l,��;������Ɉ���vq��>�z��U��ç[��!4ڰI�PW-\�c�_.�|͗j0�C>l�'�Gs<��=\u�ޣ�.�1,�i̽(	3�B�<p}�aM�Ef1��H��գ��^IߵeFGn�Q�mm�y{�e��}��	��Q�e:c>c} UQ�.���G�#�6����?�c5��V�+��=B#�;,V��!����W������g�������]��EN��o��Y�w���p�vE2��k�{�����W[�$�犝1]�rh���Q�,���J�r��X�߾E����n��L���EY�O"<S
<���Ir.E������V['��r�6R�O�h���Pbbb�^� ����
o�]Ć�$bvVr1n�(]��m��Z=�
3����}i���`ΰ�C�j����͋��b�N{Q(�K
�s/B1�T��P��%$z��B/e�?�X����V��:11�n:L�H�5�Y3�E�R�S+���b�����Hi#�l�'c�K��R,��Z�s�6�^#�a�M��x|��)9������1�ږY���c��)��㒔}^�x$���P��P�VT/޹���BVĪv�#cM������\h�]X)��2N�-( 0Q�����9ҿ�:FJ����L��/�K����̗6�}�Į��4�yI���~@�HZ��|�4Za:��Nʽ���d���S��Q���΂�����=M�vc�� U����mxx�T�zL�u�n�j<�Vw?,V�x%���o�{�0�`/n/-���O����H�b޶����5��ё��J�^\ ��z�bae��ﷂ��7�`Y,����}�1\= �я����c�ƴ��S�ȿ3�4c����	v�^ �lNQ�Ns���������ֵH�3�{�#V�^�s��KD�4r�˖�+F��dS��^Lv��'v]�tE?��}}�N���B1X�Y�!� Y���ܵI	&�7g��(L!�bi'��O�5/� �����������ߓ����H��0��<a�!3�6�2���O����f4�9����o�n�ł��?̭.��}|���z5xV뙼�r�ݫwe�A?�P%ְ���5��U�֧j�?�u�a���"���/�V����R&�@��a´5���.
Ë&��	��q�����/S{d�����i�;���*:a�*�RSnO"bR��A���.FD"�^1�	����%�9d�[5�2�N%I�XΔ���꬟\"��A��qD[�_M4JH�8�r?i	@ç{��*��44eX��%�?�,�Y���u0�w>��=��l�t	Gǿ��t���<��0K�ܖ���e,NNNN3�� �����1hդ	�����x@�=�h�Q��^� 3��9������Le-�b���dɣ������+�㯆7Y^��J�<��S$��<{�v�'&8�a���5F�/��)�z�Jk�	K� m�>�l��#N$%�hl��Ldy/Bh>���k��q><�q�>��Żrע�0�*\ގ$��ϟI����S� Gpr���Ab��:�+�TEcb�|�L��.��px�~4ZE���$·��p�Veg\`/�9�+��LH�= �얆�c.���-��RÜ��BB̮���,�\h�m��dU�;-��ފ{��z�_C �+�N�������z�S�/�q�_���W�z�$��kk�g�����ɺ���-�|�qO<�U>E+~���J�"e�EM5]s'*y��e��}��X�b���_ʁ~I�
�w���~S�H��P�R�����ms�{������=�N�)K$�&���`_��\��)��1!�ʡ�g�9��nEփB�y�>�(Ǚh�buۨ�4�v�?����p��H�_j��Q,�w޴BX������VT�m-���I�4�`��[�:#I��4�R?M�cz����4��x,��lYZ�IYf֪���/R�pP���Ts�!''�V����b�5IH��HH��	��G��X���5��@i�y�i�0�-��/�2�l�����Y�\O�Uy+�>�%�����b#O�����s��3
=�.n6<\����(���yqAMM�.$�V#��R�ҽ�ڢ��:}H� l�"\����ӹz����>F�����k\DT?Xlbl���)�,}�TS�x��F���ɂ��==T���y�s^Y��0��"��XP�}���Z�"��I������%�=1��OZJZqz��+ދ�M��;N���4m8��gb���v�Es���<�y����JM�*������}��$l-��2d��-{����?�o���Z$������:�8k  $|;[cǕ}d������\~}�����z�.�Ub�Tط�Xȸ�B��np��IKC����Q�i��i�Q����w��a\,����sx���.Fk~~~o��u+5� ��76M��k�7ؕ�kU��F�L���Z���naA5�M���>6w�.�|a����T�E���YcY}�hFAA�2SCa���Sd��y�$B<���ِ$�����Ͽ�V����L����f�dH��z���v�'�".{��0�l\�k+��3��f�Y���\#(<�.���o�T�qy"c�M
�@E;tj/��A�c��F%qIɌ����͏t����.���e!C���6�z��0��1s����p�F��j\SV5�7�q{ğ{����{��3��8X�?��{���Φ�Q�X7b"K���IQ�0`O�^LL��זz�H/*�?5��v"�Dr����w��[io�[�Tfaaa^��G�W�E�}o��"!H�H��)��t�"]�]� ��J7�HHw.�t��F����Ê�ĝ{O<�9�١��ԄB�uQ.B(��:���ب�$`vJ��P��4�j���9�?n���6=G��JѦj������6��>��2�i�؎��B�^��V�90��#��������mp�җ	^��)-5��$�"�w'���d��dύ�VE�^ �1ۺM��BZ�A����*�����7xb��B6[�2�E"�Q���`R9M����Cztaj(8pu�}ѧ��n�esw ��~̦��3[2�T��,2x��GQ`�.���_�,/��g3ݣĿ\5�,�!�q�<��QiڼT������H�J+&��始�m9
�V��R&��?1�)���sV{�j��H���������9���uJ��'9���''�b`y�[[|<!XIxsu���xw%���Pgh^KP_���DxAv-����b)�C�͜���a�L����^j�&d:��ʵRGBn+��j������T����.g;���� �Y���\M�=><,<��>�_�[�E��JRؘt�6�I}l-��Z1����a�h@�������t�=��١SCC�a��|/����ߔ��YЧf�k�w�l�KhP[�_��{���s�
������yZm P�%��㲀k��.���g@g�~�AQ��	��v��p��u.n�:����g��m���r�+�i�u�,")�Y0N_'l T|��m�x��=@8�
 g����
ri���_���XTP��h�L*�>�jBG�K�f��ƾ
0m]��+p��{��/��C�g#�,s�����C���(��H�Đ�����d�vBΔ���_��S����]��	QIXQjް�X�ť�m�P�7$"�����a�4H�a�%���؃�L4E�^c��	{�K���!B����f�˩��s�BJ��"��vɸ�n��3JȰPĝ6���$y�J��$��p����T���}���u�Sa7}1�-Q�_./D��#ZQ��Q��Ā%��l�}�������=o��eڞ��kB(�;8��J^�����	��A �EX$��A���5~⵽x� ��z���O���E�4H����f�tHM]��|�	��w���LN���V��Bc�{��r�̟�&S�'��o����ڝ�P]I2��2aE|����ك��C�C�&?���v�R��6Ln�_$���m�d���㎍���ʝ"i�I.W�<X<�,/�r�)�� ����R�Bʚ:$$z�_���d����MO�z�����S��^����	/o�����s%�%���Tҡ￵#�^>��n$Ż߭�׌MWSI�J!D�!0�/9��!�֭Lh�>H�/��/�q��Yᶭ��̼���c�yz2����g�X9��c�%تƨ�-vEE��NE�7��ԬO�(N���/;�/<e��� jX(X(���¬����P�����Fvv�̙?G�{���������j����H�,�;��_c��id&������&s)yD����x���B��BG��/�k��Y/���������p{�y��3�4~u�c8z���|1p���b;8��|�7/��q��n:|{33�MO��^�#p�~,����j,`@�CB���L�̘�D�n9��D\>E�I�{(�\�Hn�3�ج�s�tU�Rvuʹ��|1r�J��|��$�{�x�4����]\W�=9��[��s�"��6���f�B�	�k��AV�$�@4���Tl�<��i�W̇����-W $���:b�[@�2���F�RLQ^\R���$ϴ�4�x���猅�����|�X,����>�U�yw�Y�W�W�moF��f���
&�L?20K
Z_ �P�ܳ�<�MO�����)�M\gp+FG.�����5�l���~$02+Z�q�]������"��!��GJ5��t��̗{�o�������}��ς%���W��ŃL�߹�#������+�Q��"T7��«�ϛ� �H�˲@��	Oe��8j}��EV63����F�����iL�������L�՟����Q=8>鵨���ߢ}քM�ģj{Yg��1����DO����v�lE_��-��U+RD_ƴ���7����
��) �3�i��j\�� ?�0M.�A��ְd�ݎ߰�.��zf殭˵�hP�ܾ(]�0��!dR��D���kC֖��P�6�i�R�y.�Otq�F��+�E��~���٬�3iJ\'���#���B��8�L���|S��"FPGJY�+Q�s0C�C���7�d�vx:e�RqS�
�c�_�y���$_��y` l���6�[!�nb���R����44*Q�"#�aZ$ ]+�z�+a��Te��1(�*�?�>�.�4��7D�~�2���N/��gVҭ޷�O]��7u�\���m��c/���J��.�c�V���;�c�K�M��=x��ӓs��I����>��x[@@�W R��|����0�q�Ԝ�����	��_�]�/�� lי�z[� V.�'�Wk�]ͪM�B3 ��Tedxx^�bU���.�%nN���������'ȅB�b��O����W�"Yxb�_��e뵽�`��[D�QkD�f����т�¦�τ��]J&*!�?���� �!Y�;�)M�sV�j�99kl���U��;�0z�,4yd�mO���7��
Cv��R>���������Ԕ(�7�7_&&�3�C�4����X�����4���Tz��������U�c��7O�&��r��?n~�����} �Pe4�s��Mh���	�旎���G.I����҄���6��}cx ��
0��:�SۧX�g�N﹫S����T��
��LfHP�a �j0N������;mmE{�T�gC"o��؆��LT����%_�r ��A(Q��ٌ��r���`OxI	��y3Ri�Xc.��H�VwO&�9�=��+�z�z�(
�I���D���Nc �w�d�ݶB�.�a����2�e��`�y,B������dd�����i]'?���A��*߻s}y��;7,H|^\z�R��|u ��'�kH8�=C�NF�Ls�֌$�؃B���B��P'�@a�s(ڢ�'P��P�1�t���d��������|��˯_W=��ݽ�m�GN�\�#<gggO`
v��rX��wg�~��)�]����\��}�/��-���#��J�o*m��!��34�r6�E������oc0�cl�r���9�D;�:�S�41��Z2`*���r׸������iB8y�I�!ѐ�P�s-�(� ���]'�����^�����Ql��r�R5Rxk��ej�������G}y����}o�|)l�&*�@/����.��85 ���tq�/�ظ1�*r>�G�!���1`����^���~v�\�M$U�]�lX86	�YW)�f'g����y�����
p�4Z/��vt?�Y�k��B��,���m��!��3���{��p�"(�	2��Ϟ-�*��)�g�b$�HZ����B4�^K�:G�PR�w��葤�2���:)�5�%��Lk���1C@���
�p��,4�u�}`g'3���(�.;��o{E��'P-��9�4�����щXQW�)0#�!h�cV(
(N��!���L0�s
��C^MՎw�=qr4aX��{�q8.4������<���	$�TYM��Q1Q�9���B̇�b|�T��F}�I�i��B�����~�E�pAN.CX�/!Iϩ.f��_i˳���8��ȾB�x�@A"H=��F�j�\�ȡ�ѡ	@W��z��J`4�`Ա���-
��q�ݍa���h������O������#<�)U�ZT^���o�����_�ٹ�XL�^N�C-�D)�`@V!�T�f!���P���zmqc|2��i�H��+X ��|�+��Ȼ���=�T��S90��!^TAϝ����xAoF�����~�:��4D�'sW!MB����g��I�nn|v�o+�.���D�/�ϗ<
wY�^��;����n�}��Y�]w[�~ǵ�@��˩t�\t?�-_�-;���	�,�ߝs��+�yc~"j�U�m�d�רkȾ!U�Tg���BL�<Ԓb�o�!�POT"	�w��e{z�@,3���X�W~Z�����:���s���Y�k�p�:1������`�}�e�������M"��uw�Qlsg�F7�k�F���X>������RCN��(�����V0�R���E6ǹ��DFчA.�^3q��� �%�I��Qu|#t�4���Ri?��#��!!>���� B���{��ڄu��yo��@�!.�5����e`�l/n�nc�q!z�q�a�I�s5�7I̚�}���!�Ä,)m�=$&�$!�.�E�0�H�J�VL[��)�ZM�[nV�XT��\�vT�[�c��R��Y��0�b2YC������HE��GQ?X*��U����U��x=8�v�P��tS�5ÔN���q���N�m�߬�"���D4��R#"Y�w����3��T�e
����U�B�P��Fi�P��{����j�4q"\�?m�}��y�d1�Ӯ���E�}�sOO�C��0���Fz��J�yn�ӫ��L�-��	�56�l����O��K��^�?SS۽�9���"�İ�����f��/�2��MD�6B7��j��H�����@�>H�#�q�Y%��V����U�@f|r<M>�"��`$㸜�x������U|Y���~��!��l��m'݃W�S�X�,���LK-�K��7�b�?�"1�kT�S>T�^�v�aKj��^�F�N�j������&��P.�=��te/��Q�c����I�7֭��f���Q��K�Z�</C�	}�Jr��+��z�,��-J%Z[c�4�_�0�W�Sx��}=J��!��4��	�Ē!��D:��K�~t/�gEuv{襯奊��[�&�?�)�|S���doы�p�?^��c3m�X�ީ�粏�ZKTK�+�+(��-��j�������+0�����*GEr���?�王�z��rց�Ҷ �~�aXO��mu1�&�WӄO���8��U/wixx؎^��O���f�{�}�^L�Rr���F%}ku2o��������Ĭ�JPиg T��~��	2��XF�fRv��|���V��×,���q73�W?g�����^y⟺���K~595AT[�t+fw�?�\I�|[~�3si��u'�-�znc�0��'sr��PQccJ�c��R!S���K�qb��̻�WGk��=�Me�R�	����SwHF5��_ iVp{]M �D��ȟoV������|� s3B:�e�G��x&7~�~ t�S��Ѻ��~e+����9iX�b�෣�|��T���k���ҝ%�_�UY`�!�
��Ϝ�߶�7H_P�U���٣��Dz(��n�hGă/ȼEg�	�r@N�ǯwJ�U�L��(�m�I�W�ul�Pv^�;�xQ��j�����Œ�~s�@�!>�j��0챯���i��l����5��Z��	�?����}�#���O|�㈺�h�Oc{�;�i~
�D�:E�~0���9���%��)�e�������T��mt�r�%�]3��T`���rտ��g%G��1Y�؅�L�#n��#F]�u{|;]@�wP���ˆ_���f��f&���K�'��1�
j�w���8:WdX��ע�G#j��奓O����\SQ�.Z4l)�,�~�5�S�{��BC�J5� g`i\L86�>�76&m;е�6���ކ�l1�$��-����)�nm�0�>$݇���lZ�D	��eb^_�z}xd[(G�*�.�~<5H]=�s��'ڝ��䨀
�j]fꅜ0|�2:�Y=�=x:��T�&�a/����H"W=�~L�KO�Z|qPg6=��b�x��N�,� �E���N���Z������އ�q�8���=VZޔ�*~{Ѥ.��R��Z>U��k�GJVY��ɞ#7N��O
p��=]�+�o��ϣ��5��I
66'��U7��Ogj�]���#����ত菜!C�W6�.3�Dg�_f��-t�M��Ro�/�͐������'Mnn�z\\��@9��?08��Ez2[�Rw+����8�RGfWE�{��A�Y������j����ޮI��I��\8��{�^�ˣ�W�/�����u0k����I�~��ʐ=/�v������u�3�5��),e���](��i�\ �PЋ	¥z*$�>�ѿ����5�F���vB�V�&� y��{R<�>�˭����D��n������j�D�u�,�w������q����۸��V'��sTE%�?sή�)��ƽŎ��kW�+]�gch�����=T7�<���aU�
} ��-�y�|E���t��C����>ç��zMd���Q��,���������N'fD
?��6���cߢ���V!�����e��"V��d�d}|�jŭt�V^.O�O����	�}�t:n|�k��`
�C_�յ�H�����x�[�˵��g�Z*{a��8�_ɕ��j*x�����Ѐ�g\��R��pn��$Y+���y{Y����!�%�$n���ه�TKO'�}*󔃲㢄À_z��\�����[Q��K��q������}{�1�V�2s!��:[x����@_�x{��`,Rĭ~|b9�Z�pP�\0]�p0�����G��͟�쀻[✄��)>�o͒e��;UC�[W����]w>�U�W�-�N�<_���$�,/�R�Ψ0n����]�˽j��c1�Q���s�$�&��v!��2�3�� &w�ͧtug�9��մu��Ϣ7��t�p�w��󮄫ݱ��;��G�L��A%Eh��&sPX>̨K/�Q͛�r�y����C���/.�)y���ZN��j��K9�Al<���3~�n+*�Q|{_M�~��6Y]#g����x�xo���[d�]or��]�:�p��J���攔���|�����*��i���wym�`�4�{Լ��=�䓒�+U�~f�%�|�0�jt��'�A�.�w������^���ݙǋu�X�-�_("Sl��P��Wp�|/]T�N�2|�zc^���IS�қAy��'�s�����b]�tX��o�uC�m�7�n<8�(0_�X�C��x)�E�H܍��~ݶ?�r1�_�i�>:��	���0�Ǻ^xA׻�s��Þ��������`�^��������D�r��LV�y���F�r�}@�s�c��9���\��}���=H�]D�+p�<�Q�O8��<6����9���؛��O%�
P�u�Ǧm;Y-&���9BХ����t�>媟�ʪM6��p%
�y���\��$�oz-�p[\b�V�,����:`���Ig(ׂ�
,�#[���q�deǱ��v�y{����K�8�I�X�^M�+����z�����
���+:;[�[m�z��'�����6Vp 5��\YY�����z���\]�w�P�"��x��ˮp8���x{{�ʆ�ɿ8|�=�n���e�L����ó���Ԣ�,EE�G���99��7����J�=\l���&湹�5����B�.��%_.�'�z�~~�8�i�)�Z��W �l�p�������]m�M���'�=��?9���^9�y|=ҷ+ �m�����M�Mp!C&7���.��J-��<��ś������g�����I"��5��(��2Ą��W��n�-U�����ltJ�����	�d@�� z�.�u4{��[1is�y��̮O�����_��s��9F
�/N�#o_�Uޏ�v�J:�3�.���S=��\�Z���X�bLP��bS,��G`��Ga����C����.�%��T����]
����3���oI1�}�n@�og 	���봄@Y�>�vHAX���.U�P��`DO�A��C�y�]{H�*[�%�`�÷�R�7�jE�es�S�/��n��ZϞ����!���ow�J��0���\�>|�6tԺ���ڰ�dC�d�<dn�i�Ɗ?����FLD�(WWǢ�k�'m�0����ON�z�S�\��/$*
ǡ�w�_7ʆj��	�3T������Ԍ�-���O�k���Ԣ�pR5V����l���}���^��R`���^lwz<x���9�*$W�Ü=m��s.��Ѹ!S{=�kvg�v)L�tI���p�i�d㬸��a�-�v���̓''5�ߘ�-�����-7�*s1>Á���{�ݐ3�V�4���>=�]��;*::;�n�+х�8�ˈ6�x]�X������8Ӻ�Z�zؔ�����.�sSV �r�]�|j�f���^n#�&1�m�9'������n�W��N`W],� #��)v';!�&����G�M#=[L#����g�ecH5�6��y����(��0��9��xM5� a��f��\#�^������Y��D ����Ix�v&,��g�F~�D>���ي�B�,Y���{�r_�����o�����zaXނ�Ӊj��_���ߨ���k��?���fOC��#FX&�#d���S{�U�"�-���w.JgvU�4xu���L�]��#DBܗ�<�<L����з'K���>�������=�>j�\^��p��� �'Ư���^!�`���gK�4�����"QqO�+9��}|d��
�>��<���L�k���9�~p(!u�1{k��/t+C�k��cEQ_�fߴ���E^R�g�-����Mn6c�k�-��&'��j
zN�f�NƔ(�IK2ԒA������i��B����������y���ܞ�YJ9��ϲ��d�����30����r#�Ӑ:4Q�4I1��	��w\�rY9G4��##6/PO,�;��X���Ȇ8T�L8z�>OҿNJ`0Qz@�M�ۨ�J#��߭�Lcd��X����Nw��b�s����TO,�XӜP��b�ײ3s<�h��{]�v25th�~�;�?V�W��˿��������,����	cQPB�l��Cn֟q�f�Ejv�'&��j��#� W߸6d�^�O	`1_]u���>�j>��`���׵��W��1�'�=�����7o�����U˙'������d(����`-Ł�AYplG(�Է15�S���Pn�6��@ZᱨPc�2�p�['������_��~F��ƕ}EY�H�O�� Ѧ�V�{ �֣��u��s�e��ő��T�ѫ��ٌ�.֑�م���DJ��H�t.q�هزU��!�%��T�C��&N����o�������|�ښ����wʈg���5~��[�pʩ*+�w�T�$j�	�����/��Z#ą��z����9 4H�ݢp���:?5�B��x.�rkkR�t�l�ì�}�.6��'x	��CnE�w�t���mD����x�~���D��Jd}IY
��Ȉi]��A�Ч�]��u��h�,�/~Pиz����ݱ�ʟ�����i�������C�a���8I��� �����6is%%��c�j���7����.>T7o���5彍��w�-��;�D�nܘ��\c��jl�v廿3����6�̫�X��l���D�Pe��OS��ҲX�7���C 5y=c�638�{R�d�X�w9���&��t7��|%�N�h���8(��A�g��h��>#������I(1p!��1�����Af>�Bn�K�ؔ177׮a�#�����ߛ�bWo������Y�����ϫ�8Iȳ���8����޻�VI��5�'�y��sZ� R�)#u��~����N���<�陘�5��������=G�ĪIhڙ�U�ƣz�������<>I�?"N��I��!��8t
�	J8�Sg�p�y`��N��{OCYR��]í��􎿛9�y���yϒ]sa�G�N���$0�����H^3	,9���=���܁C�)Da�Oe�=1.����֓'��?]����VJ.�;���9n߆e��,.+��|�7.��?v��ʰ�R"7��-��`w(�<E��#��>���f2�;ĥaZ��X����Ӻ��$
��^���+�q^��"74������sO��a��ל���<�={�3�,j��ʂE$!��>�}�`�9;8AK��������Rb�g\�R�&LTST��8QT����fU�5�Z��9c'L�/�YBi�$���9}pma�]�pD�q���+�nJ�!�Ռ�L��0կ�[lۈd�)� /��ԏ����ʘ{���=�|�^H+`��`���v�-s�ZZ�����y����_'���~�WCn���԰M��ʉ�1�^P�a; ������dJl���/��_��c�Vu,s��~TO�U��w�[!�R��x��\4 ��W����[��Ճl�ԧy.ߨ�pzs���9���1��@~�� ߘ��1���7�#�����+�or�m� |�#�F���"V��!+�}�s;�d����P%�U��W.��=�f����Y���#�D�W3��]:��M�_d}w�9ل�� �ΰ!;���xW�tv�t�o���x}}}�{�4�FLx둵��Mo� �	��~�%(	�>��b0�w��0�P1PCa4�4�Wш5Y���<�(g���!aU]�[�u�} b��]� �y����]�p�FZw�ʰ�����?����[�FT��}��O䈢�<P����"%_�w�@@���A��a��Q�H�c�g����B�w"�� KMo�A�����.����8�	��0BCA���`�	?����nb*4{ݑi޽PEL~o�|kx)0�ӓnn�(9�?G-�sߐ���\G***�ĕEU~m����ߝK����X_�vv=�����͈.b��i����Q?�<5}���y� #^'@���DQ҂OC� �A=��A-��J��Q	/0�q���x��]�T 3�j���\�@��Fjaii������w�( �%�cvK��8"-��b�s`��a�c/{П�#}3��&�`}J`G�����8�ofл��;*7<@�jI�8x��߲��ժE
�+c��,�u���*F��|�]4!�@r��G�P613�}�j;Ů���ս�j,���U�_w͔����Mv\��K����x׍�VOn�V�8����(V(m,�b�Z+T	��s�6�D霉l��`XW�5��&~֞nO�#q��L]7��������y�l�v�4u6�����=;8����IJN���rt���W�P�	Ѯ����~�+tmm�+o�������hL"?ܽ{�Rcк�����/�9"� ��:.e�5�H#�Ї���:}y��
�b���T�X�(��_�D����:9��˭ |�ߛ����|�3S�uS�[�g8�Rr#I���"�A�.D.`�F{|Y��D,r��Mr�����АȀĐ@� �mږ@"=P.�>�7��9��/���?�d�b�P3�A̑������ވ���H�i�2��Z�"�/�0ˏ�؅�k�̼M�����P�.�OC3h|�1�����D�(��f����
Q�02 d�s�Ϡ&���A� 2��f&IGd�)�C��n�9�!���$��%$�{��]@� ��|�g�
�FܕF���;}�Ŏ;j)j4��Ͳ0�4�'K�>ڡ+�.<�]x���c���J�`��u |���*��4������u���u��!|��S/��%¹4������I�6�3V��m3I>�QZ1�-�'KLmP�]l�A��x�'_�xo��N�I�*�����q�Sq���2U��ъA��)[$cFx�j��&\��c_ٝ�B;��5gG�}� hF6��9Q��:��q}�]�uXs=�.Bk���bv�3�#-�����l�ycy��珔ΰ��3��q/�y�����^<�$	
�N�m�No���_�k���]WW�}Қ��/9O?�7Ki��}���u^�!<�V[�!������*��:�u�'6\s������bG"Od{Y��mP.��N��{�
+]gQqԬ��(�$�Ab��(��gs�jCbAT��`�KKk��H]���Դy��c5����:;�����5�<�[�VRd㲹Z/+�ZP��l	��}�e}���F�:��i�*΅�ξʟ�+qF��é1��㘕>�9%#!ȕi��k�[RĘ=��z��U�N,.��S��]�Gw7%�0i<� أo�G��62��6�,�[�<�2��ї���C�9Ȣ�/c3�κ�U���+��7$�Q;���ܛ�K���3������&�Q���v�ַ&����ҦcL�����|þ$� ��u?���`A
5�gο�E�b�;�~{���|C����C�_�bK�~��y-�Y2����/0ڼ�q�8W�u�ճ:4����6��8�����k�(�����&f��X��&o�mS�b�3�9!�Ht�Ky$
2j�f����t]��/(��/d��Gs�~������n�'�Z�奒M&7�-BX��R˰����X~��}�
���J��R�`�E�����L|ӯ�9�ݦ��%,��J8Gg ���~J9^v�<��MP'�'9:N'�,d$>����W��������̞���ě���X�и�Bf|����-�j�o?���FdɝO't�D�a0�x�#,���*�
�i!�����	)#1ј�.����fH��� �P�������d��Z5K�\�f���[�2�o'`SrT�N�&��%�*&z�nl��6c6���J���e�y��)�x�$����4��?T�#�j���qJ�ؖ��&|/'z?N|F�<@JL�G����ոЫ�����8�G����<�ң�[�[?�YE���J"���Ȟ���.Rs���݋�7���~v�""�LT�Wi���9s	�yպ(������&��bs��;�������;���֖��~)0 ɖ{�B�r����aS҉������RM��YR�Ύ�Mu"A��JTS��>8ӷ���g%�t�,ENl�IK
�5��zմt�[�$�{l�vDv�jH��f���S`I�*M�ů)g�i!�l�� +��饢��U��DB�R���Ê[� .p����o���^5�mw��-|���ƨ�J�~����šu*�Յ�����N���[��A,��cs���8�`��f�l��a�&�8��]��A���fz�<�_��R;&��'^��'j���[�1n|k][^Y	�5���%qV�I
&7	��� ��t7�a��l���kM$��D)��xeuKK��tw�h]_����w�P	�}�g�����9�!J��Y���ٖs_��=�`�'������;Ӄ�����������[�[���e}�ud��r:z�}�Օy{�O@p�[�	@H���y��8��_Ç̅_��Ժک�X�_�LE������s�b��sr*%u)2=�������n���MK�S��QQ� ��=YjX���uy�?�Mq��ͺZ�ʜ��Z������LWb�Q:>�g��/ȥt4�I�P�"�|L㈣�u�J�q����d���LNSru�ZN�����r�6�d=c#�E�Z���+��'fT,���5�f���N�^x�[�g�b9�P�ק��M{x2����x�#q����npM��Է�ӫ��Is�~�a�\o��a������̮�<^XV;0=pJ�N�Ӧ�Q�ȣ��5�+���Ŧ�I�u����z��������%,O"j���O�v���x�ar=4���2��)Y@����1pF�g�@���U,~�T�f{Tdj�7�a��!Lݝ���Y6k{�xޚ|rX;� �5���f��2��V�v�)��9�|.��R@.�F���if����$ܽHt~�d&��]���ó���Jɥ{W,����\�H���O�}�*z(C㉄�x�%�Ǔ�A����<k�W�%6�]�T���g�44�ш��m�.@��a�v�x�.�r\Y)HT��ԫV⏀��;rV�L����^�,l�L��P#�o��'��z%A��y��[���&��c�xb�MM����P���M��m��l��fmll
���+�,�|����5t'A�nh�dll�h��������CQ��W;��>���v�U^��3���2���_Z2;�����N¿{���乾�\���=�ӝ3���%PL��c�LK�L�oO}�A*M��	�S\�X=����1t�\Ovl�ŵ��BRqY���V��eB�-!��)ۏ�8V/���o����F��	���l��TD����O��s%U2���DB��uM��7�M��W_�q��`�@c��s9�!�n;���y殚���|��]�����9�����d�����7@d��}F��0A��uy��>1���������.ۮ��y��Xl	+Z'`��3g���� �>e��T�n;%�NG[��d�n�?���Vg�[R�M9]�C�C#�r+`�\ 6�lFGG�0�i߈�M���H�9d�ٝ���5��?K���>ʤ?����p�5/`�B��Z��x���\N��x�7�T*U9���՞�!=9X��}-bo����F3Q\4w/��!�~˹���� k�y��N�c�δ������:�>g�p��[XRbX��O�Z1������ /�
˜�FJ�y���٘��o��non@��iH�7HQ(m�{(����eP�j����^�6�r߫iwװ�яI��>���Ɯ�5^�IrY@��C��U��p�;&��y9.w�(�~�-�P#���R�yz�[-�/���O�;n.������Z�����9�61Cb����wEE)`�~��
���V^j3�m�ԁm��͠*o���s����yi�Y��,W)�e�:ߒ1���L�_�:\�o�����bIB�t\��&R� ����p��������TuI���,��b�7|��G�喃�������-����X�>r��l	H�T�������
���y��c�+�P�S�\��<���V�-�K�E��9aA�ωd�%������o�bs}�pp��������kG�
�:�ڤ��1���g�����^o�9��c�a���!-��tM"�a��"ӿ�
c��MDd�v���V�t���*)~¼�
�p)���P��N`��X��8��ٓ��G�����j^���L'BX�e@�~g<>>�SmW%��ٱsZ�����"��� Wӧv[k}(��d�78������e�/�ٜ���ޜ~�~�����3m�T5x��K�Z�_ۦ�Q8e��_�upE������-��^N{oO�7����n0R��Z���Ɉz�L5�o.���ZTUR���Q�wC��a*V%��	K���&���ۿ�p	�Cg4���l ��@�Y�-�W0;R~�3ӫA�?�ǿ�t��_	��R���A8�?�Ǳ��1sh=�t0�]z	V$~�&������1�����eaG�	�3���Z;��w�>s���25�zd��v\J�q���J�˥Kj�/�I�-ɵ$} ��\pD����"۩���	v�..X �)<ɔf��0����5�y	j���Ո���aXg�<x1��>j�b�V'��D�Gw'���8��ؾ��3�l���G��$���S %Y��]��e�z���
�Ѯ�i�:`k/	�Q������k?�d���I��e__JkKIiq���q#{{ԉ���RCݹ�7�����/a�=u��E;3_��{v���:����4{��-�ei�v������f���r����а��9�`9E譴�pH�E|��~WX�xbu"���n�L�������
sż��"i�`��j�ßOݐD7G"X���_��r0���Um�f�[R���r�$�<� ��wA�g�� �l�q�>���؀{�N���t��-'k�����w�ߛn��H;�ˊK qh\�^� ��`p��	?�?�!`����@����XgK:bQ%����~Q W]�qޟ�֣\��z�nA����vt�[WX����$�P��	�b��q� #tJ��6 iE�&y/��1�A?xU�f���i�\>E��i+t/�X0D�ڴ[K�wu�`��c�����nl����4>;R����\���D@Q1�u��r�Ef�����|p�Kơ��U�n�UEcQ/{.l�Q���--u¬ǻ��f�C`"���tÂ�:Ɇ2YN��<�+n �vpY�]���6u��t��Qxn��M[K���&�oP0�a�ѯ�&�c�vϰN-nnNc�ΎOI`��s\"�Q�Oo������N����*x��,�=NI1Ϩ-zL.��찇����]�[����v���l��z����锩c��f�sN.&�Uz3��a�k-�f���]1I*��/8�w�nہU�􅜓s�l�`у+��Df�u���v��-�8�	mPPRR2(>rS��R�d�|�o[�8e�ɚ�L�T}��=�:%�j�x����͕��œ;��?F�3�`ɑ�S;���'�9��U&&�P�g]�jk�l�<_5�������	R����Q�Cb[X eU�������rx����Cj�`� �Pړ� ;N9�m�-���|�G7�������@��]Y�s���L<7��,�(,)�}�o�H�B#˗���R��a�m��%�FS�g�q~v���9�7��З1S����赵���2����]�����~#���F@�eM�;���m�8��B㏑K/3�i�~κ ��\����Kªj/v��Q�@����,��]�A�}Q`�wۭ�L�`���c���pPP,@ķ~�գ�"L��yڮc/b5��+�*��<��ds?ݚ�Y���{|6��t�M7}2��jU~�抅���fF}+z֡�o1��W=8R���]&\�["����^��XU�ϭҺz\���%��:&�)	����̴��)�u��?_K`��\�,~:Cl�4Z0'�nd�
|����vg1������\r^�v�9��K{�WW'U���
�ee��I����Qo����?tJ�tw*��) �%"��J�4��t��ҨHw7�ݼs����}�b]�]�s�����9����`��+�[g�"VV��$����>�u3e��,�+i�A�踆�����],)k��pZ�[��a����AU�qb��S���Vb}�J	�nW��q W(G�L3���xsd����ŤO���e���o���A�Dq�cˑܻQ����"���G�O��[�B?'��hYZ�n׹��P��/J�[gy3�3��1�R�\̼�����#�Bѵ;]3�kQf�ݭ�maY^0�){M������=%�̬��W��c����
xNՍ������zbBB�Zs,ō��y���89Y
���_�������K��@��c5|���L9�ݖ/��y1
'�x8yRF�k��7�'a�����F�����ǋI�dO�󣅿�r��<�*((�������B_�[�.E���L[��E��v�yֶKj--gg�tW"��+�J�xgM}}��G�%%�|o���UUW"��s��&��A��n�d/��ټ��ބP���9�ǵ8��D����Q��*��$G�+�E����6ah;���#����@_��SY��Ҕ6�ҹ�Z�`8�5T�W|үt"m��ժѫ=��a��h����������l6.����)���Ҥd��(�֣[�F����2͖6�T��.ǼO�W]{X��;zq7c�{��;I�3p�?d$��V�O��\�dT˘26�:^��E�Pl�'���I�E-S��a/���dE�n||\O-�J�)��~+���� �o���v�6A��ؔ?��E}qtMǺ#>���?C���;�:�v�uخu��w�u �隴y�סR2,�f�YYK���Ǣ%$���@R,���Y1Ap�qU��F��ZA6y���~���S`,د�4^�y����,��mօ
m<
����͉]��U�@[�"SfbR�:�>4�Z����k$��W��"'��D5�g�����r�s��]�3���#]B�Y����qB������T��T��XB�F�a�>�A�܂���|E߽��)P��n�&W:��NKj�3Vܟ�s�`ȏ�'wQ�ބV��E�ƅ�a��L�F���L�Kű�iǇ;�,�}��RQEI$_�۰����U�<�(�%J��ꏌ'�x�}
_�Yt%��CǙ�Q��Trcz/���Y��8I�#I�8�̻aƎB�����!=Ghc�]^�1j ��phMB�6�G��^�%ۢAW��l�haYo�S|�gmSQ>g��.����r���FӀ�b<�P��~?P.q�'ޛ�^�HЊ������Tj�/��9�ƒ���~��vc,x��iЮ[Wv��V��� [�:�~���[{�C2������5��@O�%�9�RiG��F��wm�iuԔ2�G[P��t<��P�� Ŵ��֮�Wa����*���$k�����Q�1�6���)H1�%6J<�}M}m�m�;#�W!,�q���}��F�Q�c�t~��c>]ڴ���D.�:J\I��ų���//|��%��a�K�>Cp&�f͉��j�)��X^l�Ǩ���&����p8E�\h3#a�N>ZŶE�922�q3�w�e����c����:A�?BX���41�Sq:���G��w������G"v��|K���l�1HDk[���J��=���e(����c�ڷ�)�I7><d){���o��!޶X�x��E��fT��ES��%n^/�˶����Hp�h��<7֓©<�-�$vB��5���h����$�~^��s@#$d��ҧ������4q�����dO��0v��j[]5��Ȗ���=���zܽ����]���&T��_�~�@,�g{�za5)e��-��aݜ	HgB���)a���k1r�0�Vk�h`]�Ϙ����=�M�(�^��U�n/F�.8�x��5i�;��OC%�B8}��c�pꗵ«��,������\�M���-yv�,L���c���UEʱE	?Sϲ~ֿ~�,��?�;33��x�M�j2�Y8�����v�3F�jo�5�{=5�֎��������\����`����U8]���;�J[&��42Y�2�s����=b��Ύ��?	S������Բ,��һ9��O����db
#rպ{hd�^d!Ò&@-�.=�iC@)G�K������\zɑ���{+�S
}q�q��v��^�sl����f�l��ʜM�`�[~9?�n��¦"�IKk-�	�eE|�V��X�yy �i%7�Tĥݥ�$W�X)C���#n*/l/�K���ҍ�l�M��Ⱦ�)��5��#6F�:<�M������%zmf�JC�3:k�:/R�au��Y�^5o|-5L9v�^������q�R�y�0X���N��5�ϴ-3�ڎΐߴ�smcb�+��&a�JE�Ћ����6,dŲ�1XJG�� �u4���G��t�%��T�G���T���	L'	ٷ��&�bۛ�K5s��T�<l�ѿ�A|`����������KQr'���7��{�_��M9mmY�'U��O����|Uj0y���|6慚�6&����*fvf�W:�&������w��Ww�������_ISH�F\���;�>��sΗ�HT{a��T��m���5g��K8��Z@��p�)� �3�⺾�3��{_3����)�)lA�K"'^n2A�����7}�+JѥN\*ާ�ZFFFc�.����o�qG�Y*�q`�'�>�:4���Bn����޾���6���f����7��������̑�e�/q��]�2���>�s�D�d��ҵr�!�/��v���K���'z��*�˵m��d?���qL[�������k�f�9����xS�%SST�p���}E�v�Ժ�#*S�C~\��N��~4)+vvy�Ҝ�;����R����nu�Ygv������9>>.2�l�-�?C�羣��i4 ��<��ո�ٸݵ
��d� >?���H�I
��a^lϵL����L�^�U�LHa�t��i�(K�f�����iP"}��W1�iJP`O���6���/\���(4���>���'��P��Y�"/a����=����,�0�r�߷�����[^_���'��KA=��kvy��!�lv�����h�����-FD[��<t�b��>���r˵���th�������V]�EW8.���
�#{�|A�������\
�u�8��uy��s�����g1��U]6�V!��͔��&ۑ�����������60P��F��� ��q����VS0��lll�~|�mo��Mt\�CG]�d;����������>>��M�F�Ɓ�m���W}3u�g[�줥��c�oG��N��`��;O��Jrs����_M��7|�F�}���l�MK �N�B��<En�N����KC�7��BKk��pތ- �3�lK�O�8����x0�����kwo�I��3%c�=�,��"s�����&�,WWSv'�C�����\�D d���{�&�+�'v�e�6c?��Oz�3ζCb+��_:�.�����@���Lp��uuu����i=!ֿۧ�˿�|�0D'[��`D�IY�<�����E �}ɍ��M�jF�> �N�
�ĭ�.���Y�f��C���|�[�nB��+n���S�/t��^�m��ŗ��hh랶��X���=�H�&��ș�eEE��^�p��-��"a$oX&y�eVe���^T�2p�1f�R���U�ı�t}}9��m_XQQ�ٯL�DiDaEl��e��-ɿ�}����,h=�k��R�ƿ��y��/{%�P��B��;̶/�����&WP5���_~�?Z�P���\���oDxaCAH�Y枯��d��N���Ԝ����C���άpU��΂�Ku\))���E*��"8^5�x����Mou�ˬM�lu�2}B�on<ʌe�Q���K+�QV��
�o�edղD# ���S�gWTp���SG�"Jy��3G��q���E2{v����=���$F�Ρ����?�g���p;a�GՅ�����_C����Iʶ�:��Yj�"�?�"8w���\P�a�A���	��C�E������������o����uR�_��`����}��Ri=D����������7����,q�H����ŀ��<_}}�OOl���$�#�³�|iii���>�>��:�z̧�ĹҾ~ݶ'Կ�i���ywS��y�pKZ��F_|Z�]s���,L�����ہ&S`}��h�1�V�q�s�V>n,Md#��q�,� *���4���D�΢�F�\~Me�:�q3���	�x/�\��j��̠-�P��ÇO���2�ɨJ��g��Ccb�A�s��\�>����O�I�:�w�L�lڲ����bQ���Q��5�Yh242���KN~W�<[���Bx���{�U>gvD����d�%:�PgEl�K������@�۷s��˻��aς�_�M��<��F"���G'O��ds(e�������&Wk�&���q�n�4�1(%=���v߱���).������~bLKuQ^�q{B��_	�h�]#(�YrG����þ�o����^x�!��/�����kTQu�����X�����7Tkv�c�"�l���2�����g���I4a`d�TƁ<]�9�m���*��5�aqlЫ�ߙ��δ 3jD�?lŧ����4���ԫN,��v��:�[�o!�BD�6�&l�a��z ;oJ]MXTu�i���m@<��:�����.���A��bf3� AX	\m�m�y���5�B�D.�_�7q7��)g��	c4�Xd�[��g��A����Q��8Ol���9~��\����f��C�����O�X�L�y����u���~��� oC���S���@�-�||u��G@X����MP�'�<��)&��Y����ȥp�h#�	E���v�'@-J.���@F���։B"@��w���I��`�F��M@K�9�a�+�K>�.�k��{��"��HZG�氂�*Y�q�A+Mx�nw�B��1�ӳ�q��o���<�77?��	���ã�~d�xBg�;4�_�c�����+X^Z
OKX�_�s����������jS�ʬ�u�����kw�u�q8r�C� /���ʝFTf���<m4�9�(9��K������"�kj����y&Uf�*��/7]���&���O�0
i�3E[��Q�[<��p���QL�=1ii�A�9�t�e:?�g��~�=��⍄�>������߉_[<JI�a@V'}B��j2rOQ�#	�ҼK��c�����������vqP��c��J�#	d��R�S���p�~g��Wrw���O���Z�~w��:t �.T)��iw�Q�>��g�:��j<������
���C�JF'1�g���u��S�	�3m�"�F�j �y��l`t�WOF���I�{.ĉ<�MSQw�_���}����)fͳ7T�^��.����	s����{�{�^T�d1��E�t�w�,Y����i���s�uX���k���`9�p��5��T��;��B�@���{*�u]���@Uk5%ߕ��pw1��7pk6�i���J4�O����,Է�Ԡa|jiNl�2��M�c��ņ�ҷu��ÓPc���NFB��ap�(���Vv1�ua��0�/*7C�k}��Aw�ֶ���+�}{�P���RPDDY��,2"BJsş�e�H�0�Z����y��u:t�ł/���)�Ϯf�//^���YUfO;���4�)G�|MnO���P9l���{/����G;؇-�_3��oO_O`���2~�ӹI-����5UEJ�j�D�Bx�H�jF{*��;��U��ǮmO�᧚��u��?c���8����H}u՛�Gq���8��R�� �p�(K�2�%9p8�H^>��}-k[����CL�p�U�����>�і����J��2U������i@�dm�������t��WG�4��,���)g�8�չֿ6��|�֋��F��NV��.�7T���6�a�@�l����;���4c�D2���KF����� ����Yn�\~�V˿[�0��5�P�[i�{SFcL� �W][�B6�(M�������s�, �3q�y������ؚ�t��[>3��`��*�>`�2�OZ��pP�P!��F�y݂����T�B}�k�~rO�H�������,�Nsj*ҌS<eq`~쯘ӹ����ͱ�.E%����6��^�F�����nJ����n��kѦ��~nG�b�煳�[5��:�ς����?3�"a��G3����� �ܕ�Z��������1P�.��Vp-� 1�uj�"��`LdAPI;~�.,(X��3Jp��~��_����/�����g,�\�f;gBެfg?�n����n�xuV����wK�D���{�"��T��H�d�xH����j���_o�$��d7�8Y��k}rƢ_[d�?[�2���@�~�c-HCE6>>|�ϓW̑�9�a�ӟMa��덶_���w��2V*1Tz�������q*�K����6������Hܫ'���O�9����!]�r��bXPo�t���k��$�6?oV�>�_++�@���7�Qm###9D7����*�1u�����gd�x_����bj�7��~���hEv��W��`�L�*��7D$h��+�/���O�X�+��5$Y2��;��h�CSrQ/���2ޫQ�P��vf�t�)_���-��� �|z��Ϥ��� {���W�&�g�&��ϑG������_C�I�t�j���V�5{$�D��;(:w��0����(N��p0+�.�%"bt��@�6�5�ì��5�|�RXŘ��W���v�~��"�A�}�@�*�������X;Y/�F#"P*fݑᑑ�$�~�O�j�~Q=y��E9��Dܯq�'|���H�q>ԞT#O��v�cH{�D��"��p����y�v#6��T������4��W�47�笰��E�{����i�{�:��3�����(���gP*M�J��@�RD"�[Z[�^�xG>�0U�亹D���G�WoK_������oI��4(�caurtҼ�c�\�w+�r[�#har�܉�W;lp���U/6��b�.i�����W�
v�׶m��z�b���k���u���5V����HH��w���fo�m���/x�F�@�&��_,��:S�ko +����\ߠ�]$i<`0W�1e�*$�y�{O�Ng�o=4�(";��S�����MSB�z��:k�7���V�&O���N���jf�"-��(�:}-VB���7��ʍ���̚����/��f�Pit�EcX��S0���4�w1$�P�wHs�'rO���ύ��
��f��)����������<涳��j�\s�J�HǏ��KV)��ի��r��S8���/�6�m�%�/���|�K���|�������[XYm�1G�������)y6��)���>j}^�I��w�g��an����|=�n���m����(�����U���D�ug�x��
���2C'�n4�' ��џ��|{�ܔ����?�:��-��u�:�x��+�3y�,��;4��EA��י`�f������肏a�֎��n��z�w}�PG,W�C6�Hrǒ���g�^�l��2���{ne������FF���Q�P�^��d�v������ϟ��%�oL���g�dHb���E`*�pE��	����n��7������DI�J8WE�WEQ1�M���%<���ᗂu?y�����������E��Fm�}�+9;��s�u���rEݭc���IP������C\������L���D��zd�2���)?��Ya�}9����teC=�Ʉ�E�&��:�����E�?\��h�O��}���lǃ����k�u���O�ҽ]18A;D1��~�]�k����/��g��؞�*sy�"u����	N$&�I--��Z��Q%W��C'�k�Y^ڋ��\X����4�`�ׂk�R�'�*�Rjj8���� qw�C��x����2��^ �:���P���b�����O�]�n
���@�|.�h�������]ŧ�?�/A������Z�ھ�@Gxk&�&��<r�}Kv�&_�A�\}��}I?}���[3�ܛ�@��YuA�z2��.^�|G��t�'P�s'כ�JQ� �_L��y�@ �󘟅�gG�/�OK����0Mc�Sa�����EK�X�hX�G��~G1`���VW�X����h��ʢ�tw�z(+�%�����N�|�2�.P��O����Nb�}��1W����,N���0�=���Jx	��!Խ{��N��?*_���<0�\X����=dt��22>�4�y,89-��&���K[<��"�1��}�x�\�vJ���K���-^<.b��԰:�q�4Z�B�r�߯l�J׭��կ�G��(p���O�4�&���Jd� ��y��S����Ig8.����n��������ԋ/*����ƽ;c�)�<�y-B""�Ps��憅M�R]\�P7~��E�g�,��Cw���0����ZJ����3666���I]5�o�f�$����J�u��4=�+�.x�BkЪ�?--ڛ�����5�_.!��8.��}��#w��g*�'k��Ǯ�`2�#q�����Ԡ>��#�z1��$Q�7��~�����~jT���}����e���w���!Q�ʞh6%����kml����������[�G?$  <�:�5_�����D"Ҩ4���0���lY��G�X�0�|nu9d�F�u�D֗����ޔ%�6*mb�a��'��iw�^�,��]֛KII	���j�[o�zs��_Sm�"Y����^চ��rC�p�ˑ.�0͈GLA��ف���>����}��\��OO_��;���HYnSRRbh����Ftn��X(��Z��C#�Ⱥ�Q�su=�l���~�����&�s������`��v���Ӓd�������dPh����r��ެ����r�u��%��Ar�li�{7�oA���	�ǣ����8����ii���\ώ�0b�oy���:!k�a�K|�" ��"��V�y%uE��������hDs?3�����V�9����������'''לg�߰I�� ��ɾ��e����������j*e=V�=s�a?I	����g�Ԏ��$�2�%F����1T,ө0��fқ_]]�*%��(ࢢ�j�Q}�|�F��ST�v�{Ԍ�|������N#�X8ɬ��7ZI��t�3G
�W�V�'���QQ���%ODHh��^_��3�y��M��?�:��9��N̅L/�`��5=U��f�} v
�a�F�;���%���vur�$,�(�L�O�����8G�@�����͖��1��}^����3���\Www�����A���d�[b-b�<��Wo�������˧����K�U7����5�.F�/x�+OU��.��]z�,$.�N�E޽T�;�\���p����I�:����eZ�x�Q�����ϳ��~���b��q�\��N�APP���1������E�wD������c���f��I�Ǖ(�sX�-GW&0�~ZlO�g����D�int6?=X\�_5�.�9�/K����Mٕ����bt���:܊n����\�[Plz�IJa����+�Q^��4����"W9��N3hĨ���;]ǒA����e�e�Ҫ�D�hWʧC�{tQ7���R��YG�#"!����}BV�_�4�r�c�k"���Z��Gߋ�VV�v=�z����
��G�}$����K�WP3�*�!���'�0%
��Mq���	�e�'����mnP�x���nJ�ƪsvv��d�H�;ʠ���.��G�=��������NtLO�BS|�"N�F캕��ד�"�j�a��'�09,��NU!��{��}�����	��4�,MS|�}�5���fG�~HP	,Z)��x�C9�G���ι�0pKI�zx� "�ƿJ���C�0 ��?���6#tbg������P���l?��ԝ𤣣�����:��?�oU	�)(( -g��B
��wE�///�x��ҾE�#�HRBz�\+���J��L��j��&�����a�2���G�̨2�:���	3�r��HH�I7��yP"�E����=���^)��p=�D�^\�>	.j_����nVVV4�
3��Y��]��ɵ\R����<�ш��FF��_!���sq��V6��`d/?{*�V!d�]�Kֶ�l��x���t�~o��)y���/���E
�:��p.�	\�:9����`�G<�M��ߛ]��l���njJ�3�RD 7psàw�H9N�xyH�X�G/��s�y�2vщ�Й�W�Im��ye#e��v@!� !�mt����h�q�9<>~ff�׽�8�Vߋû���ݲ'���F퍡0>a5�ggT�o��J\`�H�F�U�/ '���z���U�����#Rp$5�|�ހ�"_���x��;��Z�@�'r�F�ֹ$R��Ky{��PX_:�U�~q�<!���򼽐vT�©S}H����� ����g|��ɬ�Y��u4�i�z]�Pp�2
	�C��;�V��P�Ԑ�à^�m��c�(J���7f�9�� !I��0��ǳ�j
caaA�}y���1@�K���������)�yot7�����ȣ�w�b�h��F�"wHe�eH��\�X`�p�O��3��r����Hp�x�	Ne�/|�4�N�X����%�����_�[�.zQ�u}��ip��d���`hh�E����PU����*1�ap=G?�%�I����|�E4�.�,�yg�՗�,#0
�����Il'���zL��Z����0��F��������X���)Y#Y�۫g��R25_;;5�)C�s�Β|�ߞ���"��ܶ#��3�m7��N��JJ��'��T�)\��냖i��J���HD9�'�������wO�X����������٫�����h�w���Qd��u��I�������������U߿x�������} &?3�i���<���"��'xoy;�A{r�A����s�b��yL�pe�OiO?_���1�&s=��ߙ�>���nn2'���{��y�ұ(��yy��0��E"_:{xȁ����m�<��<-m^Gנ~���G��kޠ	�W2��f��'2:�P��_.�q"�}�����G'!ߍ\z+ѱ��[�j�Q��
n�6>;,�P{"�F�3���ŉ ��iF�b%dT�
,�tn���\�F>2��\� v�.���A��L�9���=G�	����aǢ�q=���Ԭ濺R-�4귏�t���V��t�K����奎�/��T���@͞-�����m3!�}�2Z�^P �j#{$	�iA�|�vp�QY��w= I����2,�\^ABgg��b��0Qn�X�X�HUtt���=^Z_�<jJHH��6{<nt�K�����S$P��?�����������cr�:��lg\�@�0�qW���V�&���-�����η(��6�����{�t}>Y��M Y�����XEmZǜ�n�Y��:�<�.�=vd?E������7�!P<@��7>����Ch~~��F�Ǐ��(8��aPa=ܞ�Hm���n^f<˕L��t	[�2���k�.n3���a����Ui\E�����fD��v�Fn,�=27fe1
mڦ.,�4E8�)�#���8�
��x/�lq��߃N�:2ǅ.�I�{������2��6/����|3u��&��>�H�:Hbӭ�zT��w�"�e�v�"�7^�R�3��X��:.R��H�r�o������������ɬ��H�"��&�1(��0�_<�RH�RȂ$�(������(b!�s��H�b M*��th��ɪ]u�+F���$H���L}H9y��OO�C�MgjmS�_�Lo(((t>ܘ�5e�?+�4lW'躁�;C�-pyj��$Olp|.��$O�uG� �0���K.�r|��������� �d���:Y`�Do�B�d>U*nv�.D� �\*�9���,EI4�F���7��	�W�
�W��6]�����WW�q2�J(�I�h+�K�+������Y��31��q3�ް���:d.v˳���T�"q��@/@�V�-�]���kv�Cs�ҹ�Iˌ����S���a���J*W���%��.�Y򑹙��!О趶�Vi?tAx�P{>>~G'o�a|��V����G�e ~�9��E�5��#)//�d���dY��|5�[8^����i�y�yM�����|��$恠��D۶����!@�#�7�]��Ѽ���:uZ��=�0�$��U��18GȦ�hiL���a4���·��S[qƳe��Q�eq�؀����ך���DA�k��]��$��o
$'�_K�; �¬_�L)���IP�oރYC0�8��𫽙����X??�W�,����0IC�V{���<�H�h����$�0�v^?=\�N�4��'Z����/4Vw�A") �ky8���_���;i�eI�彼{H4d؃�a���x��w�p"�J��K��pR8p�c���1��X�s6���#��j���b]��7
	�D��Y���o0<��"�l�fg���*���6'

JkE=�۶INNN�3g�l�c4t��Mܸ7��Hvcw��f"i:UxIG�{,�TI"�q�Ж��+7����'V��Z����EBZ_TH{�>���a�7��1��Pqm�eK��5��n�|.4��͵ ��p�9��Tsd�Gd�z���ķ@�@��;���P�I|��KBKG4�������j��z��sS~�%����{x�G��0-8u4IY�=�囥5r�;lV'����>�߳ƀt���WY���^����n}K�i�n��g1�����7�B��hi�Іkܸ&BcJ ������9dJYm`4��l���H��P~x\=������)�������� X"i�399���j��Q����M�iȼ�
�B������u�LϳL�:u�=8��L�A^*���`��N�V���s���<��$�^��z�2$)��Oq��8�\Z����`�ϯ.~��O��������#B@M6Sq�����Ճ�< �f"�����ho4ml��b��	E1nhh���i �U�A��pwQM��&������X����*��$2�;��k}�6O>��h�6哅!yB_���O�_ۑ��~i��D7�Mz�!}r1���N�0 	g��t�f��H�h����1A�2����CE�5:��11� �Q_> r��ٻ�w������r�	��8����]�0eX������0A���>�犙:�B���_���n�n�m���Lws�g�	T ����oߝ�̺q��?,-�vuw���/�)����T�Ի���-�.S�m'��[��*��𓒒��!�v����r�5z�0G��Wz�
6����{�x��m9u��PQs����tU�Z^O�],ZW�O(��37o��������hΎ-�km����Я��+]^����]��zR_�n绾��s�LKL��D,YYZ��������Z��F��0��jK�f�zk���W�����w�&�=O�N>�������!��Z.� ��ޔ+J9���/�V	���:o��L�\��(�
�<���񺒒As�������P�����
���T�_3l���$pԅ��>�����<22���r!͊G>{�Ϟ�C����Jw�F�3$��Ń<ʝbQ��F8���0*�K� �d~z�G9z��tk��2C��NJ嵌��鋦��7�H�C�{��q�S:	IĠn��IU?=�>��o��T�<�s�G��B��JJ&4�����5KơFM ��u�MU�B ��`P���I6���		�������b�~�y)?��
C���U���en�@����nk�<1�˯Z����������� �!hhhl�ԕ�/L�@��A�y�.���+j	������|���r�f�i��F'�}T�| Q���v�y�����vvG3(Y5[e}R�ݰ���י���j���j��dd,Ԉ��pI:�`l�����30I!������ѧ^M>bȒO����a����������K�_8i�Sg�'ˍ��9��q���v�	z쒬��.�q����fB�P�͏V�O�������C��|o���?���~Y�碿���� W{���#VLU� �$kjJ�Տ�q�K��qĻ����h��XJ��ǀz���������4��8h�K/��U�����rJ���������M�J�AU,�17���۔��d��J�m������ �<�Yw�z{��߿��I窛�稞���,�!#�l���ӭ2#���#�;�	"��̠��0�o�MB	H̵����WO�?�3����8j�\��@BP�ԑy�i��'����9���v\M�QPV�~�E�t��9�}x��n�m�3��d�Gh��588X0�^�;dZZ�WGɼ��AX�BM@�C=�ף������9�i���TJf���TUU�5�, �u����N3k�D��B& ױ�����Z}D�>%,..������x��D~�D�=['O��oG'��: ��J�<  `k�*�2� ����o�o �4�����6�<�t������H�������ɜ�f�|h���p68�C���/���N���x�Y2���9���Zk3�w�}EE��jWO�
����X�A͞dI�h�WU�́��<�4aP�X|B���|/��z��?��������WC��
�rssmF>�A}���qp��JX��/WAA�+�/���3�Ӥɞ�ne Yڝ��KNN�:���(��Lr8O�'����("����<�(`���r�QT�DILս&��@�( Ҥ_#_T��L�= ����}m��!���-�w�T�@�+(�qX��۳x�Җ���Eď�w�_�gszb��hv����}��j�L2&�Tp��ݚ!�׏�#�����.�6������2P\5�-�X��L(��׷��^�((���
����>��_�2�N��Y.1��Ј�{{��=h��U�E�����:;˰:^���40b|��@"��oQ��c�|a������~�A^3{v�+��TP�{ �of�D"����&+L&���n.Q���M}sg�w��z;��K�A)Qp�p{` =#��b��T�56�#����e1�L��hr�@��F�l��,Ѷ�k�����.D���]�aP��O���y��/c�y뇑��T�9�} �����Ik�/���o�����\�cǞ�P���	:���%!!є��Ԭ��>P��݁r����|�0��V8\\\�fO@H�JJ�P���/-u����m���I��3���۟^��t4�J������%��N@`^ކ a�m���. -�jQ��*@-�'9-�^Ւ���T����u�Q���!۫���i���� Y��
����R��X��h��&Rr�Z����ϧ��/ K��d��>a�8u�������Ư���(� �=vÁޣ���&�f���\�~ܟ���w6���4�]n�R��bjI.S¬�3G������A;�73OB߿�.��W �����W�U���}��r�wk4�I���(�����*ω��.+�n�"��`��d��i�yj���ד.~��s:���[u�
��pě�Lj��>=�-������_��BuB��~b���� D��E�@�h�Q��sx�?e��O��&{#~�/V�/������>}����tqu��T;X�X��s��iuO������	Ȳ&s�}@�^G����-��g��D�0u�$��A�T���p�N�mQ1�Ӡ���M ȸ�������!?q��/��r��{I�
 ���g2�����g��_�>T;BKn*���zF����ǆJk(�~W�y�j�{�p�����r��NذK H���/#2	�b�؟�ȓ�����.�;��hP��G�TTTh��p��A�Ïd�����^���� �r�}M�ˌ[��U�w��"?Ro��kt��ٯ�K�g��0����o��q?�>4�}a�'�])���>��/oG담�B�I�P퉂F
��wO���!:8�<2�@ʇ�μ�ʸ���e����ɞ(��}���.�]t�6pVr��'����Ƌ\Y<��Ҡ�?��Ǯ@I���Wc�,%�{��_�	�6�I_�M�V:7^�i.����Hܕ��i	��N���q�Y1(� �����\��,��h����_�noo�o��~ Y�I�}���yO��ɟ/���? ��hƞ�����ɽ����[����,�d'6�ߞr}�"���͟[���/���E�[5����]��!�
D��D�A���� ��	
� ��
Q�L��������Z�F���|/y��?9���}o2�QIx�B56϶G{����̠- ���D}�1ٴK�w� ������ �����K���Ҭ�(�w��d^qy6�o����߹��o�p`�n����a?�m�;#���î�\�S5��Zl����6��ڐ��gB�@�%��VG�}�q��(�� y�#q`	��2���-�f�m�Wx'v<5��l�*��22V��+���=��1�8 dٍ�E��.��7y{\usq -��oe���7x���k~{�\1�c��n���߽���@̑%�f�#[�Z�W������wj�cM�I?^!!#��^���H�xD TmG1;��)kϛ�h䱑��οP�C{�5�y�#ƭ>�6~gFA�s���VId>:�� ����H�4jlS��V �~��I�����a�L�w�����O�'�U&"9�������p�ʎ-��ԍ��I>{�´J���w�_�>t*����]n�	8.��P�Uz�l��֨�IJ®/Ud�]�:��#�/Y	���_O�?�������3n����EF���xi&�Qi�7�d���D�p��]�/b����;�ҥp��Idp���>��<��>�i�ϱYY�qt�+�فr@"�7��%2�hֱ}���ʊ�Q%5�5=��&
VW�y����X��r2{����f�Ud�����ܼ�K�t�%�`hh	�쉍�a2fPII�ZH,���o��d�CY��h��?��:�����V�K��F@	�K@B�C�2�Q�nE@���A����w����^��B��}�Μ9gvf��Y�``@;�w�.m���;'�q�:D��_~�9pڗ+M��u^�u�� ��B��c=`����^TU����:�B��γ���͝������������KV����V�q����n8H����p�E%�=%U$Q�u��M�<JP~\��T)�����ў4ϳ2ի��?����=� ��R�K!���+A�vS%�Bbb"����H��,|m�˗^���y��&��4�Ep��2�GL/k��=�(���FL�up�����g�B}}}�ӆ�~/?���C=M�c�<�`0���n�Kă��)>%e(pP��@i7~}��*1������_�[[[�>�~ϵ�E�k��f�����RL����/w6�ү*���o�t�P���_��;��8^�s$��%v����4a�ܪ���k�|B>���_���WՂeVQ�S�8���nn��b�e��Dg���O�HA8�/��LL��I!h_��~���@��ִ�W�aUT5uɴ&> [�G�z�Dɇ��_� ێ�hQ�\Q�J�����D����q�"���Y� �q���@B�m灪��`������[28��xo����=���,Ѭ���;_un�P	[얛���O�ư�3@QQQ� `��<����,~-2؜�*�*}��h0��mҵ:Izn��w2�-�M'�˴�1l�סr�+b@0��J^$Ʉ#�: ������F��i���bu-�����q�4l
���7��j|��<j�2i��y'�]�,,,��g��NJ�����W�o�{WZ�!V P�p�cgWZ���t3A�(�g�x.�FƑk�$�bY��n��c~�<̘��*��t��|�}o̲!����Y8#�!��	:�E�*8�e�7��$�����"/�6�'7�43V椰~E���o�3���/[y�Lઌ���s�>��xme��q�1�V#� tr�(����$��N�Q)f)�9��^���"�cg�͚ˑģgg���~Sx��1�E�1�����H��1
���!%��d$�8�y��K���jX���9���y#y2�!�
KJI�]���,
w��` �B���g������}M�#h�OS����E|���4�"ý,|ml�	�N)ݻUD&s�!�-���\f���	�i#�"��Ϭ�;�~�G��p�ϭ�������V�
��.��8��H1

��%QA��74T�<�RgQI��'���>]*�Ui�l��?�s����^��{���o�T�;�t�ܭ�l-��˾�+88��b��q��zSJ�p�\h�-|��_����T�E,R�3k�ߛF�=ŧ��p�}3F>�Y�:��f�� E�8���)/�v�0{^�J��ɿ����|�����M��/gQ��piIuu"�!��쫚@��7~�:r	�)C���22(� �K&��!���$�Z[�,) m�
��� M�����8�&�@[GGԆr�������Y$�����:\׵U�����>�Lb/�/����~Vk %����73e��GH+ň�g7�$�^#x$��e��������B����"O� ��� ʭ�?b�<M�%:�W�cܛ,(<c+gd��.�iI$��DM1׻>�D��Վ_]��:Zb�큲L��H6��~���KC��~�\�/*i�#�*>�(��
Q�7Cx"�����"�2��o�Gϭy� ��!�i�jf����qss#gpuw���	��B���זĝ�I�8I� �Ҫ�ҀE�D�Q��55���7̟����_ur�g���SX��!]K�=�?�,1��Y$(�R닩�=>�鼪����&ȉ3��[4��/���}X/)�%��x����gc%[�t��))�i��mƘݩשD��#�������>�bɵ�v�=�ToA�N����X��3����Z�O�����by�:66��eRRR�9� f��Qqi����/Zڸ茁f�6n����{�YTΓ���r�LOw�yE�dj9�?���e���)�A9JLnmNI�����J���ra��6ky��ʠ���0�CAI�铍����ȷ,9���$\텮N��5m����|d����V�(�#�0껹;u�Q�q�B�w6��6fYO��ے?�]XZz���d���\�_�&3:�[��6�1Q�I�}^����:�c3M�ϭ�����*Zۧj^_^̣F����R�c!K�W�2�����,���aoA�%�1s^������lH��r�4���SW#v�#��zb�Pn�%�i�fSެI˖�6+"��s����]y���Y!��-���1���[�߿/y��>9y܊�F���W�����W��`+� ����o��P*ĲK=x�F%��Bqm�:����a������A	M�G���?D�%�t��x�{������7�Lx�v.@0(-`����>�=�#���iE�E��Q���F ��\F��|��3���⏕KzK h� ���P|��ԃ��l��8bbb�oR.��߼yS:��w�)w�ȵ�ׯ_�-���KW��.p���f9�)H���gx7ޥ����t:�m���MF���S��#F�Q��"��T������<��3�)�+��gr���q�)l���`��΂��Įl���K�G�����c�C�bH+��N�;,(��W�6@�!���I�Ӳ�Mu|�Kޟ��8ϟꆆ��9:��r1�����664\U����-��`�d [���$8�%
$*~�O�-sZy��q+��י7�hU<�k}{�x�h+�(?i����=��6���;W�*���Y��qs��D�Qͫ�0��=kA�]3�^��4k~#�t �����?�����E��+�p �L�7���OxS�=hw*��~�V�������y�|Tp�X��[�@�>2��������z)�?�3=���0�B)F Ѫv�#��0�D~x�N��?�!
4�9|a�-fCI���/��?�]�9XL
��Տ�ܕx�V��F���?U{�F����mV�v��',�ӟ����4��������P�m���7��_�
�ۖ}W �=���WA�<�����9�ח����6H���m����s�Onl�<�?0�&:���X��h���B��4��z%Z�V�Ĭ}�ff�o9m����7N�7*�S>���@p���l�j�|�9�~;7v�>{�B`�z)|������j�[
~�**���H��Rg�}�oV�+������)k��L�]!̆�U����q%�w{�y�$��S��Ƀ���9��~�C�M�T��E:`.�����|�}��C�݌��h1���J�ן2E �7��I�YM��k���?=�8EV�uz��(|�m��p�~j; ���w]p��O��PS�+T��ɀM������M���T�����/-���ۛX�����.H�_$^}e��φ�Z�4�"���d�^�>~��/7��y5�ԃ|�۪˽Z9�.��O-�q�[�X���g���r�����h[&���p�6�ҿ��uNE��ٯ=c��I{$D����QQH�������..��'[M��ȯ�AL�����;����q�#�G_W�p8 ����T캈�gU���1�c߾�dh8��b����~�����s���{yzw ��3�`cc�����]�n���066�qa��!4m9�sCG<�0�G�F2��yԫ]���>���ړ���7?�wq�94s�����o����&���ϯ�^��Cyr���H�!��Ɋ��>� }�Ј�?~&���y�
y�U�X���?���6G��x��s]�$$�檦������ݸ������IJܭ��G|67m_.|��ߚ	�{�����Z��ǦD_\O?U�>���K|�*|�e�}y���n�3GZ/���8C}�m�j;Q��|���x���"6�ո	��K�.�T���A�6��տ~�'�>n�R:���_XS����T����I��IhJ��T�刦'_��Ud������L��R���.(ڿ�_Ss%ʅ��������ꃭ��77ˁ��q\|0C���ٟ=Qh�)..N�����<�tEE`�����:�gri;���Ыjh��D�m�H�3����qc.[w=ڤ}Q6��O\=.-����=��{�1��"���$y�/K/�,-��m�k
������z����#ﴴ�$�J�R�u��Eખ��N����:P$3 ��a��'���
��L���R�\���_�|ٿ���/_� �m����X Y��>xs4G���W"
��U}dM_h�����35��zk��y:V����7�s��~���SCjb��A���-I����T�5����-���t�'^�q�S�H�?꾚��(h�v&"���i�=�!K%���ȘH��s�Ā����3h4�ҡ?�?&>���/�H�G�ɄS���I�����j}��!��d�����<|:�kܓ(��m{�#�hu�@U��]�֖�ho�5�,&'��@��?hv��GE��g���*�����gG��i3�p�����:.�w�0	����=��v	����Btׇ��t�,�O������ZJdHg���Xb]}���aa!���w\�U�^��2��}CC%�v�>{v#�5�P�
�����qZ����6.�qr��1��d"Ŋ�w��I�v�llfVJn��Xkƾ=�\\^N�r��ZD�0X�s]L�a��V���6	�P���C?�[���9����.Nٗ��#���p���f��p��w��u��<�v�Jl�/kS�F1*���F��1�0ȗ��>�I����wX�M�("�I�.�ݕ*:�����#MC,@�����rqQL���q��įd�@�����<dŏ���xc�"F������|��@�x�ӄ�Qb���tww�=�XVv���)��䞿ePNZYYy�kna��/--���0�1������&"���>;;;�\IZr�pʐ���bbgQ�,=����ˊ�Ƕ���
>*L~��:VJn%��wQ�o��*����^���g]�y�
}��jk�Q������/4F�#���VL>x�D��6�H� �՜35hDU�oٴkE�-��uK��I��&�E��î��MY$7��E�2�C�h�=��=�D��@FBB�c�#i9��N{�bo�tK¥[�����m�S��<4=+kG��>�A�ֈ1�x�{o�>��i�h
�
{��Mb����D�po~~�� P�FCq.b^�'#��S���ޝ��G|�(�WޕD�i��۵k׮\��Y,�����m&]2)-�_���@>��*C7V��|O'���©�
Q�A��������O<�،o��l�V��aY�à���54r+"���Q��n�`n�8�H,y'j�ђ a��F���Ma��O^%��t~y�e��y���1#+�-��{I%�\�z�=Y�+����	o[q�#���G'�<(L<�m�~�i���� js��f�t ##{'`�XmW���}���a���΢^��T��A�$�_���D��?܍�_fg����Iή�5���qPbl����x��r�I�m1tŻ{D�N�Rt��b9M�v\������ �'�|��E@�iӈb����gs��\��yl����Lrt�2~�K�D��\BQ֍���|��H(�c�W	/]Y�&'|�'=���m�&K�l�-"٘���e�5�*��B0�J�[�b�,ocQ.at�ƙ��Cq���A�'�idp�����)�K��odcþ�y�...�mg^�W^Jr򅚚Z�*;[�qqq�2O-#?����<���I�Q%0W������y��W�����imkC}B��?4��_�A)W������yx#���~���2���#.B�b�?/�~U�t�ͱ$x`=q1Ek�����e0���ϭ߱������hi9���WO��1�7�J-��!i	�]mR0K)j3^���\䥕�u̝)�3Ma����7�W�wEEUV��)�����ĂI���*��YeKK�0�������\6pXYY_.��젢�D�~mN�+Ɨb�i|�cvC��'��M>���5)�������&eg�vM��nR[%ֻ���Z�� O�_�+�7a```ea�2/!ONN���`qѢ��o��ϣݗQQ�u��yŌs��)b\Q�D�@>~>��7�R� 3 <�c�.W2��S��&&Ҧ��]�A&��}��,S]����l�󱙁~�%����	Wu�>�%
�ޭh�{��ܡ�Z��D�T�MRB�y��A} 0��)�ظq377����=q���m� �r%���}p�4Dң����_N��e�f��{��|F�(���ީ���E܏��v0�a���`.`�=I2�^�x4�{��X*O(p.766��jHh���֭[�WVΟ���KHJRs���wp8{�	33�=��ޟ?Y�o*x��M���n�R^z���(���7y?�q��F��+�Rb�}�WTD�3J�������czc/����u���ނ���LE�ц���}IKӜq��&ak�/�U���;�7�BvK��Մ��fP�=���/��?�wvw�|�[��Ξqss��̇���:����!X�xK�Ͽ���MIƏ#�E�NH�H�o��3�^�����&�\�ؙvw��O��c(((`�gƔ�^vuu����rY�V1+L���555}��(ң���?_C�=S�ݝ��T������3��������'�0��K #{f> �h�۷o���_��J͝>�z��걝,oh D􌌴7ob�PE=1��ԤULvv7��!	U���P��]��)+�	�0�R5��yF���l���x�AP���^4�0=��}G���k���Z:|�e6tf]`ڔ��{�XXXP���p�L6�3c���u�᠞v������AJ�H%v3O�F}�m�2�7�p�  ��O*`�Eke���G���L5�Y��bQ��M���`aQ�Q�)��BC M�b���陙�aAק��Pq�j���������oD�P`nh|T
E����N�y�[Ab�Rrr		��[h�-_GgI�a���5I�9i�D^��g��݇��k:;q���_�U����;���k�%�=b�3�иϱ5�BX��D'*Jegg��Gc��&%� z�&� ��i{�N�"+��ʓ`aM1c.�r��?2�L��滻�x�.���6B�����=�r���z��W!�傺����Vr\'�5Ұ���g�e��E[̀�0���N��藵_b����mXe0Y
���+00ؚ��BW�sJ%'��P�o;3P��`a����p�@%��$�h�>��������؛,~w���߷�B��'A¿uL���o3�` �!!!FO۪܋��)@�涧	{���o�S1�L'���n�wTB�ŵ|�*/O!�����m��6)==�Ĥ��ɚ󒒒�q�Ѷmm[r�Tw�._���u�㵴��^�0T������O]��uy��7��>]��[[j��!�7�䋰c���n޺�h���@� @��9b� D��'�d�gIW�(=�XPPP�F666V�����_/R|����D�&}�қ�؄�j���Bՙ��唆�=~�+����9Y*���2!�Ҭ�`����ND"�ğ��p�9.���\+-��O�{���9���חyy�涾~�v�<���&meee�D&N��0X�_P 6Q�957w�����ip%���� ��rF��L��94����͔�>K�`9��b��>�Q�����������%��b9�66���q#���U����j��mek���'��MI������;���>S����{��*ܿ��]��32�"������K�����ZB^'%ս_�<y�r$��T����_��U>}��1>wf����T��������U���5n^L�
�eT}�y��sxs����/:Ntݙ�HG?{
������K��W7��G�8r��99����w��%"&���=K!�N����<���/b1���ED(��-�V=��ˎ
�탲�gF�V��!N-.2(��1ޙ����1(̴|IFH�N��R*�[�w0]v��f#�i��	��ʜ]m���7wv^:���w^��>;��7##C5xg�E���Sg�S�#^������j^�T�桚A ���z욝��e�����$���j��;�]"��r'�����zwm���Z-ʪ��:,��m�P�>�7���,l�՞?���@fg�^.�~�ʌ"¶��&#�>�N�q' q�{�L��>�ʃ��f�5��m���Qz@\��x=R��Y�Y�����5h F����B�?'�k�Z����m��x�]��_�: #�hh��[���z/_�ٛ���=^�H������/L�b������D��h`}��Zf>###��q$��^FDD�ש��.�0�a �i98��i@��f<KO��l�5,xq')���_�O��R)�_.��h���4��HE��6��鸅K-���b���gjhk�;,���𡙢�"`�3�P�`�B�ƶ����Ր�!���[��BC}��x����
��T>��T��{��a
�'?����T�eT������a䤤�[3M��P��(�	��(�*�$鄧��,�g|�<���Nm\6��h���>K*���j��66b��E��<���qd��IHfNwP1J��D�.�knf������0	U�xV֬��k���G�O|�[X�������_����#��W/��4��ǋ�$�$s�[ll�@�,W���s_��Ke���;�E켤�T�ȈΪ���<Q��?�b&�����o�^��>���q�NN9�4y��h��.Vv���������\���)�#,GGG��g�>�Hܻwfoc�kϷ�~�l	kgI"���@ *��q�_O1���������,ͼiXS$*��a�K�"�a=���+��G�K��g'�^��yko���@���҂�s$x��6��踞<}:�����q�e},C�ř�����G6���C�C���=o�o��F.�~��������$��ayy1��Ô��z��n��ߘh�@����H�u0H��x����`�x�Z��ub��+�jwc�H
��-|}%%T�w���Aj|ꟗ�]D]}��-|����Q�����ߊ晕�,4�2�;&}�&eW�㥪������S���6�^��1A�����d�>����
B @t��p �����*++��|���OiI��p�9�C�yr@u4�gR��(��I𓍂8������e�&Dȏ?|�`�N�Mq�e�*EJm�^��ʤ�_����)pqqѨ7Yu��687���Zq333���[�aÛ��00��������y���?礢��n�Cꡪ�+Ӧ0��5T�������,,�����j��hi�2�㺻!���� ���=Xݝ�J�f�����`����9]7�fgg��z��J쒪��e�ߜk#�����lj%w6]�!HM�ưbI1�yzz��e:�A�b��^! DvPn�xVdd�χ��֫��2���7�ꞎ��מU��$��7ʗ����v��EH��Sx�=v4hEzFF�A�s����,###�92��nK�ɉ�� F�V_�A��U`V\�G�lڅ�����S ���⪪��H`�˶�>/������2%��������,plD��G��{{M&��=���/dk��3l���i��������Tlhh@%�8Ԣ!iʟ��7�U�PF�q�0��i��\kAl���mm
��%||r�XX^EEE��
�rs��y�U���� \q��u<���$!v��KW�'�u�|�u�}oߕ���R�yvt�'��0>>nϡ����]�g`]`�`��+�(5͞ 6F�pvX�111�tu���C"�e��;zѻ���m��m�����%tD7��6盟���&5u8*�l1��b	�J盥��ڨ�������s�v�C\�������4���o��|<�'On�Ӡ�5 ��/_��k��Ҥ*�1Ɣ��'H\����\(p�P�ӥ`G�KK7;���ҙ�p���j�ٚ�����l���)�h�����?�������r�͇>�=ͷ����Cy�	�{�~	��yS�̌^O__�� ���<۠��6J�tH�X�Cw	�?�=�z�Kttthv���s~Q��Bg<��+ݥ���ϰ���Q�ďx���ϲ]ä��	d�\t���c:���ۤy�����A��p�8�kP�r����o�ϒ��ֶZ�Ͽ%E����O���n�j�6hL��r��;�Dt��]{#��eK�"���]��T �|i99����W�����l�q4�a���x��y{]�~=���&$�B<f�  gü?Y�siooϤ*���w7DE+G��y{�{��xw��[�Ǝ�0(���R��斖� `�>����S�X��CO������ĮWr��=S@�$�|�B:������e��c�X`�Mߞ�]�Q�������eD����899�� iAg�(��ZE������~�$����@i:T� ⰹ���	�7�a�2Ǜ�����q?��?�> �kXC�H��-Wt$�oTs���
0c�KSm�-��Hk}}C#��?�̓Gy�X_!���t��AgLL��R⾟+����+���NO�~va�H;����5w-����8%*压#���0�^��s��wW��p�Q�:���cf��Wa�Q�l���ֶ6��F��/#��2xX����yxx�)V
'�*B0�4�ߢ�����sNz���]��]���j�1o%BS�9�P�/��M4����4n\�v3�~
V�h�(j��96�X�m	b555��^����v��#�L��V��`n�oGu`݊��k�+�D��<���c�UUU��Y�iV5��6~b�/�a/aaa��v�z��/0H?z�ڷ�4�<�K�<�Np�5�vƶ����μ"Z4���H}=�~__����9CCC�{1�#���Q�V�Y���Њ$�:��޳���	
B����9Vbw���K���'w��0J �o�E ����Z���<^l=�V��ohl��윷�i�Y&����t�?����0?~��k^4�(^��Ū:�O�&�\C:�^0(����0�,)XRR©Q����	qu���<\ !w��W��V�h��װ?S�������DH�񋉎���B��v�zB���F��1H���F��˵Q�^�sT����!R�vW@��B�۷IP�ﳪ?��������"6`(AƆ��
>���WR����KX�+f��x���`��sHU��n1 �O=n333\O�$edX�k�Ԝ"䋴����Ӭ϶TOz!g���~��׏���v�qՁH�7L�r��Y!x�xd�靕�~��U ���Bg���7�_d�zhZ*�����&���HX&�{��K������QK$�y�Q��?ρm�^���0/�&��p;d�������ⲥ��fY��5S	ͅ����qط�l�X�����\XhODs�����fffq/1�^��(]�"���ݸ?�����Cd�uk��!�E��<CjԾZY)�}� ������ ���/X�@���[�n�����QxBPT�ى�N���m��ڵi�YW01%�̒{�^/�j���!8�~����'!q�����r�ζ�0ʒ����<�$��b�11�o���@O��Bl��?.JO_��HP[[�j�"��n��5>x�������Q��d4�A�q�M;�R�0)�b͐,u�����>}��u��%%�,�N_U庥e��bhh�*��M�{�*�l�ޢ)%��#���Cڅ��[�_��K���&o.f*&vUN��p��P%���#苏�-+kk|"�BBB� �$��W�h��yZ�cb+bԓ>R$�bWwda����-�S27���.��Ue��A>ʛ�e��d��g@�,0m2�{r�_\��q}z��`8���=�,�O��mI�/_~9�"���5�A�BkC��,�e`�!��YMe�K���F��OyДR��NJ7 x?�� �5�����0���� ֞_X�)��[RRrv�_�+8x����8�6��Z�Tll�*s������T��9J��9���	S)�v0�f����p^ˇh��,�Ο���=~�p��k�kZl��T��ח1�O�7�L�+�	��)t�2�1 @V��gt�)���������eְ��W#XS�u�r���g�sr����aw9aa����w�z��qt`4J�%�(H��m�
x[\�v�8��F`��	���ͼK��@�PPihU��p�1j�G=ҽ?^�#9��������·�)S^.�\��Lf�����r�����]?�\��k�!2-Fz�P�"?��R��������%� �,�EAIY𨃬��,H����d�2���0�伦��69��IDw��b�,�� bV���D��5������$?�h�k����$��ȐUT|��@|��%4�Db2�7��?����������Zg'0\���Pv!Y���)[(�
�ŏ��`�­��/~����:ۖ������z5�������s�:�)�����SRnf뼫k���7i�2J%G~x�]�:b�#�Is�y�gY�@�ǝ/���B:�bc�ѭX�=I!��O�A��[�y��@���5�!����an��)b���4̙�º�H���^Uv�	���X�ͮ���7��{v���׎|{����xh*��ͯ�۔��G��	P�z%���׋O ���<�;eyq�:����ŕ^M�k�qL��#eom���+�:n����Lc/�TQ��+RRR��p
�/JNZ7����Vƀ��ytx#�QR�Ϥ�8�Lch�3���24�hm�ɢ���2��q����x��V���	�ʣ|�gWpd
�ݺ:��ǀ!yrig���������5��u�F2(U7<�P���C��1�1\��0�O777�ݸ�>�{&��BΫ�a�B�r_o?9�C�������Q�]��o�tҺ&h�~�v��17��]����ֶ'E������/4L^!E���_>�n�}��;x�88�8{0�����Ώ���U'�@>`�D'���B)����<���ئ@��f��3Q  ӻ�ޕ����=%������A����WT����p��mW7�����[�W����?�������6G�t��i	bH~��+/_�����Q�/���K�yc�����ֽL{8�3�3L-
\|�g?�x��M��x������(����4�U����sZ(�cG����4N�r�L����kX��W��.�f�T%��ZÕt_:1�4�}X�E~|�����_����m���1����i�l���c7�D"if�gZss3:!�������|��6B,**�FvL]�-��n�m���̓z!����u5A���Pm ��&*
%'I��jGFP��m�o"�@7_ ��0�rMQQ�M�]�l&*##�q�Q�k{�����{~�Wdzzzs{N�����moLOW�dd`HHHhik' �D��O�ۍ�B��h����rf��,4v�����za�EA8��//SiݖX����>��l9�>�W���ߙc�d�w�z���󭪺��I�zFd$���L8�F�I��?uLi��u�b��U�"���P�Ґ��D��O��.��XnV��:̀ 7?�zC����� )L�F��k�}��KIK3���C����z�pj��Q�8�J+(X: ��m:�y�miʟ�F���a�%KLJ���"ja���D a~{k�&W��wY�@'V����Bc����O¿��b��-�$�{c�Z&�ʷ���#vƾ���MBI	�J��P�Uqee������NT=���%5��}�)Z���0�CEn�Bβ_��2}o>�m�D��%�ƪN�<�`�0����x� 3;�i�Lr"�gPA��ɉ�!m[����}����m���tu��n?�\X`��L�~�_�r�-a����\o�s�d�����7�^�$��$���]����>�6]�/��/F1��㾻���'��o�|c�5�h���� ���t����g�)11�V��E�	�骣����E�ØAAA�;��_��ޜ2@���i�?e���%;x�	�&gg�7d��,�9K)M�K%\�9U������d�I*���*�֧�O��8cHV�|wO�dW�uw���;�k9[��*z�A3�kޛ���d�lפCH_��~�:��)�2.��bwJ2�;��/�
�o���X_���E�|���}�P��mT�vr��T<�[ѽ��J�5U��W4�3F]>��Lx�w�#g��q�t�<ĸ�;�}8��[\�� 	M 
.S�y|����
6v���34��NE[K~f����?5����������O	����Jz�����5���`ev��/Y�"##���u�����;�u����:1+��U]ߏ�s�7wv��) k����P��ݓ��Z)���'�oJ��С�Ĭ���^b��� a5��^�OA���TF�kSI���?���TdA�m��˷plW{��bB"�~�~Ƨ��� 1Q|�[	h�lh��tokF�B oc"ւ�A�]�1�zee%���+��7���� h��5f �׆pr;)�����Jްq\�{�zn7"��H͖��]�y��M��)�.�!N�t|ڳ���h� .����I�l�K�`k�6���ddd�FGGg@-4�{�7���T"�9�8�6Am�I�4��<3��쫙gP�ښ�jGNN^8b���p�aB�ut@l2i��h�S �҄��>�i���Z�P���W��d)9a*\�8�7#L�Z;���#��v��eP-��]���E�Qbh�7����
��d�E[�:�8�Mf2\�/��j<Q�0�Z��1*L�s��4�̈́'�w��-%%��*���̫W9-���Qo8A!�K���}�p2�9y$̈́b��m=��#��(��vׇq�5B|�����R�����{dO8�ϴ*6M���C֢��
j���?�*�69��������]_��V�+s�)E��fy���(���Mr ��0,�:�t�,�����5�	�ͺ���7���1|�j���� k:<8�dUSS���@������AKK4�'�]Y]S]�u����LN��/�F�4�K9���fz�gً�9����Q2��D�Z��+agǁ?Z��y4�L�$9�>-��ffO����j��;�G����3i+�BJL|���D�~�_SYY��t��Ӊ�eU�����9Fz$�2��������	3<��(bO���=}8����%]SYf����k����H�����9��ЙI�8P=>N�Ɍ���\Of��O���2#���õ'C%p���ա��Fw
a�7C(�51�1e{p$!��7���{��3�6�:���K��kdM`��CyU[��Q}N%�:���%<��������C��ۖ������ �q)T ���j�����OG�N�**DNNN|l��:��		�Y%����N����%��F ��9��)Y�e��m�Q� :�6*�,vW���IL�=����򯖖�C\�S��M��q������tsx́��WQ
i$����.z������4֚���Yzy���M�!}"�@\��74�w���x�=����'՛�b�� ��>�i��	�;��l}cc�ׯD###��.��:����>K�Ȣa+zF�ڱ��V;`�zU^��o��m�u��G��6�\��^�N8?qloe�V���c���k5��Y�������D����䷯����	��qh���{zzd����ܔ�PPT�n�E���B���+	�I`��a��;��Aq�ӅGr?/�އGDD߳r+�j����.aF���i���'ە��!]����[Z�*��ڵ���$9�3h ��:�*��Q�"��bM������ "@]/\�\7:��*x Ƽ�襮�����W֣�&q��_����Oԅ�n�����A5��|�E���ߟ��W��8�;?�F�ge�vuu5u'H��^�l
%�
4�]��[`�H4��M��{:����y�@r"7��OQ����9�ـ��w����8؞����΢�|��+��;^�e����y��Q�w��|I�2�xQR!g�I]33z���Y3A鴱!+���C�\�kf�mO>{#Zu��E�o����]\\>��_,0�B�����Fh_�g�4���?v�+nM�#�8�+w��~�C���&��4�IDí���?�vc��������~/�IWě7��m���T�;�~o�Ď��>T)W�������E.
��h�Ѓ��gbbg!��/^�WoA�ʌ�_�4!�������Cb�Ӷ��^WUUU��bc�����glL͙w7�4�s����ܽ�=�1�����	���gV��� �pVF?�j
��Y��y����E��55I*��~���N%�P_/�柬���A�d�֎������x�"y?��4�x��T�t�
���#��|��`*��߈��q*M�4��nu������+���w�е�=��*��++�$G�TJ�c���.:� �|��Z����S���[��UJH֍p0r?TQy��l�WK}��ۻ�c��q�5�ULLԁr9���C�'O!��`l*Ĳ'<����w��ѓ���j
�eq����i�^�9�}Xx\�0�#�I�=�Q��ð��Cc�K]�W��޿��I�������� �h���3���a2�EK�OE��!����Fo���xf?t�1Vb�o��U�-�:�).��ܸ�f+%�r�Ԏ��Ê�՚qpp�8��?!���[=��kScO�N�����PS�g���Aݦd|�>�ādk��\p@gV�*яe<�$�	/r���J�`���.��cds�{%(�<���FQC"~~1�_���:�X����89::�ᣎ+��[>�,@�*SSN���~�~���c��t�O�ϳ(5�P껕�����������虘L���ih���>�mб6����Jr����e��900�����|�7�r�g�f����{{���|{U{���������
��� -���\Zaaa���\��#�6��+۲��ƆbV�����,-L�b5l�K�I�x���y��Ŋ@t�Hȋg*7�%�|?[��M妦�}�r����vھ�`ʟ�{Ih��o�2#ld�浃G�+Le;�B鏧���t�/&����n�Ǐ%%%�Su�&�L��h⣗�W�t�z&U�X���c�۷�I��������h�T��,�W�ɡ�
�*�o�;9�ӻ\�H@KR��p�%)�n����0{Znn�\�Pے�yaa8��a�Y���~Y���c*z�d��P1���9TVƸ�����]^�jm]>UX~>g�f���p6���HA�D�;���8:�{0������� ���O�nɏg��U�+T��L��u�>S��)��W�!d[�/ie��?w�\��-���)q��GEË�����=�qf��|���Y�7�,z����kjj�c�� ��(E� i�`����/(xOI�o �)�׫��;.S�SԹ[mh8?h/A~�������z���IO_��`E��5:�Q�[{.6�599y@]&��ˌ�|�_q��0a����D�%!���������k�zIҡ�[��)&�9���T�t���W�,�a�}��!Yˠd��;1���)	���Pr�%'��6��SSS���N���C�v/J�"�۪��km�w� 9�Ru�1�%��T,,>���͚�.\��usj����E�삫a�,�s�?����ѵ��G�����B,l�d�7��JugȎU��9�899��Wx$�/jQ�{�����W���R�c�ymmmN~�\;V��5|�9-GGޏ?���xD��U�jY�����k�1)@�k�t��.2��:`���Yw�D�r�8~l��n��nJJ8�T V���^{o/�v�=h/l�������|�hZ$$Σi衡�:�mB�rՍ�Q���u���ubna��޶��E�m./;�m�\[lL�A�WN��U�#�����Dn!�:���������@����32��hi��r�\��1Hx0���s��]�EDD�־n��Ł<C���(������3Xν�1^�с]\��u?�OFW1C�]sI�_�p�>��T�ju7Q{��Y�FEE�b�a�<����l�b�4}eXV��5 ��݂ �Ҋ��Hww�tw� �"JHK�twJww�s�����u���>3{���y������QQQ�X��|��NF ��6�,D.	U6f��>����(	vOL�*�a���sd�S$��዗H
/��?>>�	A����-�v
����7uC�����] 0����v�6#ccb���T(gf�888�&�������"Q�~�@4���.9�k��2?�����6��|4��Kõu��͏e�+P~B��҂C̮Sc5K35�Ħ��v���̭���g&��F(�����w���:���KB��I�� �0W���.P	J@���e�u��	(�\xY�X_��0�~��<�z-2~�ܹ=��a{{���4�"ᕪ����{Ә�ǣ��Ҋ+�������>Q��oc�|0�6<�i:����������>���e�J-����X4��5�o����pph�{�Ǌ1̓򲷎݈�[��F���͇�c�!���?���\.F��jo@����t�F�[ծ����1�-#���n�g[��67��1��0���D��~���ѡ~�}��YF��1����jWv+0�rLSjb�L��B�zf��'�y\�L�hm�)**R�E�y$���H��啛��솉�����m ������d�*�}}'@r�_��B��->`��N8�S3����B�K��7\��B ɝ�����Z>2r�o��22�MMM��VV��ϟ?�䙿�����bK�	z �:�ƠB���<�2kgu���	��m������爴ڧ�#��b	�� */����_�7�pq�FGG�����g"��'� ������j���L�4[ZR�V���)���,��:�����8��h����l*�p*cT�o��Y8�|Y%�;cy�lG@ۓ�D�n��^d:88��N1�XYY��P-XD�6?=z4_}����� ��M�AJJ
�4u���h5��xx���"�F�8���=k������\P�߫)�c����Ǔv�T_(��Hs�Bp��S)��hv�� 3�ȃ|��T�z���:J����QXKK����-pTB��@��Y�U�{��z�b�M���&���!���&�g�RD��H§��^�Q`���lu�yL���v']l��ת�������^X�gk8+G6m�6msk�HB@�C�ʊ�6x�X�0�m~��:? m�E �8�{N����pp`��>]Mi��  �ٍr%0^ O	�:����/Կ ��m1�S;虘�S�A�����?����%3&�����l@'�,��gW�PC]� ����V�"*���5�+|au�9FJJ^S�H�c�R獉�ASTT�D���`hP
���<�C�G�������^`݄L�6�KX�O���w�>k��nZNxsM~� �rxMi]�9�]Udl���AA���JQ�Yh%P�%d����4�����l�N���z�W��}����ek�����t �e2��!���) ����������5==}�xr.�r��3�1:5ico`7}% �=�c�MI���xQ�$�|�݄aia�^�;�;�B��qs�������fC�ڵ�d�_cC��n`�������(�����D|�*Y2ef��4D��Ղ��wX�Y%i_"�:�
��q~đ���n]�@u��f�T�H���
5o�?I��h	�SY�����z�V�#X����d�_�u�Ѕnll����pE3�NJ�(6�_ ظИ���Z� �:���H4������GKCs���ʎ��âV�w�	%*:��������H�삂�J�����7�E ��l�41l7�N�$�&�&:�AQG�ֹ;��x�7S��]� �KK-]�ꥇ�P���@�E��9�2�ZY�z�88Q�:_jq��ŞN^d >>>�lJu[XO���	�=�wt�D$$��V��u\-��@�wm��I]�]��H�Ci�g� �4cE�Ϸ5z���t���/���h��X�LMU7f #:��'�]}%�i5�W�q�Ϲ��!DH�d�����o��<��&:%9�������a�aMM���Lx!�	a&��F7G�dvؼ��ȥ,��S~�_�� ��Bf�O{Nd<<��A�)^��}uuIE��	�,�.�{��9o�9}M.(!x�G&���-   �3p�Z�QVR�$d�Ǖͯi@Σտ��u�L~�abe�06����"4�#H��#t\�OL�*,,�b]KlQ5,z��K�&����auGf��>����ϸR�m�<���\��ܜ{zr��H��Rm���v$��t�e��'ECç����emuu�`�p�Z�ɟ����vs<�>:cv�
�� ��&�-č��V�=Y�O���?5v��S��(g���G�O5�\�צ3"�"��C"�h�z��\��q9�À�Y����_���^	�z�=�'�CH�j}��Z2-{��k+�z�}"6�?�t
���B���1@}�C]�޽8)�m��Y��xqzj����ׯoz{��!L��gY@��?<�le�8���e�}KK�?T��ca(��c'�Q3]MU�
t�'ӭwx�Ȧ[���[����:�AQZ�	^���d���-h�0�i�SW2f]!

�m'��X��֥��Vx�<<a�<a���/X�zi	Ү��.|B��Cn��S�L+���}59�fQ��ު�<m������.3'��6/����gj|jd墯0<���9-��;��e�X�#��|˞���*��������l��/�	S�U]��&ca���Qӕ`�r[��k�ޯ�+�kO,0�03����-���N�3��|,9���|��Y�=i�u�*O`��޻51>��������=J.<+�s�`��s��wYYt��_��XZZ��U�1C9;��̒$������n�r�o\]�����` l���,oG�o�%۪���_��~�L.��{^Ѥ������-Ԡv�å���-�k��F��IR�;������Z���_hki͑�z��+���P��V�˜U'�]H�~|Sg�A�X���}� ���9x8�7���j�ŃB0)��p?��v���7�����2��y�iO~���ە��P�V�{3ZPcm�ȩ���\'�LD<����W�D�TYK�H�o��e8U�o�_�G�Eyɓ׺��G5��+�끘����I�׿ɿ�@���0���S�B�l���"P��\���BHg�q��F�$��Gq�O���l�JR�zV�
�t���z���GD�d\�� 6�&��2���N���9/����-u�0�w�A���s� �ճ�������zb
���nidee��ϟ?���=�߳t"��.�e�����l��r����p���׀�*N��5O����`]W�˗��X��iZ,wA ����69ʤXXP���J[��N-#��23�(��W�I������:�A����wE��Y�"�*(dW�#�͢:�Rv������x��;qq8�g3VäQ����ǟ�K,�z_��/..��M�Y"��?�����ǫ��5����	_�d�lweE�ap�K�ؾ����D�`?��A��qn���B��#������[�QP�` �Kq��G�������<v
29�SK�p����G)a3,,�\�u5>k}v��iOj��&d2W@8K���j��C����7��^����n^ίY�~����)���5Ս!�x܋��ӬAS�|6dX���~�AmZQY9:�>l8�#����m��2S��)�DyM��������p�U��٩�R/2�l;NM%�~t̺�Hnm��7�ܼ�P÷:M(�8#cQ�%����Tu�����:~����o���%�"�P	�5~�E@�0/�um]��Z���0��a��>�N�`aa}��\�A�"���g����������k���EťIBCl���w��*<��'2�`���(7I6ڷEy���l��&p���~�?��C��k�zǔ` B����b�LRW�����ڻL��H������ƨ@��	��f�5�	F"�������e#BQ��,���������я����r�E�6\|�W�MOe����z��5+b���A1�.?���Hbt�[��o�pI�l~��|-(����-o�=��� 	_������I�UH���Ҵ��`�/�v�[r��Yk�<�HH��3������	d��������/�W�(���p�*A��ۋ���zGD��ɳ�l)��!�v�Pz�B���á��Fc�`Kn١賝�'r��֒K7,��I����dLRQ�|'�y��bb��09��u4��s���yA�i�bM猌��'��.��?^|[Fc��K�
�l��k<����# ��WWW��:�ߠ?���(�n�����}��p3���z�?�ԱRX��X{3
���|~�b����{ܕ�,����z��tsp%��~�;��2>���I��{��ɩ�]f�|_ZMV{���W!���=�����U�y��F�����ihG���333/����Y͔o����о~]7H���+!��BY�]H�m[oɦ�����2��]0Z�d�i��6	I8����
 ��ֺ��5��j��L��H� ���B��L�S͆/��Mm��m^t��F���b��773[9��'7!S�`�z�����Fg4?��Ͱ��琙���
���RlR���j�7��|b�
KJh��� �Q� 	�x��3D�/K�%�r|_C����Jh�h����"�'�S��Iӆ�D�����3��7�Qs|f�S�/ss�~��y>�q�v��U�~c��� u�:A:z� ds��p�k7gP�����9���5.�"��~�H��k�Ʀ/4BZ��كԘc�M��''Z�,���S.%���9J�?TM�Y���5ӏ?~ʮW��&�������Ԅ����z�&�}����fۼ|�ʮ^��υ��������y؇��-$,,L�*�jy��?���̘�����p?>��m����0���*�$�;���؃/?
��iM�3Ko􍌌Bf��Y�x����>G�Á��SRR^������SDFFF��2H��Q���b&xDDZ��ߢ��ݡQQ���ġ{��5�7dX_�4ج�����iB��v�{�K�+*���e; F
\���6�&v��-��F[K�%/r��y$����Fu�����Z�Ǘca+v��R�
��9=/D�����6up�lM̒��ڮ����3c����j�����8��L����₊�̬���C���6�Wc��T<C%`���ޟĦh��������� G.��E��EA{���	2w���%�u�����[����� 9�{V⻠���
bgqIɿ��0��:)�B|		�������H���3��k�xE�ݗ�.,,,�}�ee�BBB�,9�l����|�[�%�����߿w3`�����<XV>�%+�}�AY��_c���K^W�μ6�͋y ��GtAY����{�cc�!�h��"����A��̬p쾨��{�Hq^��?�؇�+�0����G�Ź����c�;�d���a�����b��;aDQE�z"����r?��?��,_���iI����y�P� $���AY�#	�Ͻ��BN����ӫ�$\�)9�Z.&&&vӡt��j�CJ�$i���U��)�x�I֖��`���'o���(E������K�)��ϫʿ�S�R��y}����Jidzj�ӰF���ybzz-�o	� �)Ɋ��mP	��ޞ������T	��n 0���mm�y�y���<Z~���͕��w��'�l��0�\z�cc)�F��J�A�8�N�������}�wp���'O%$D��x�2:2�����H�F�
)p	���/M|��g�\���5g7B��s��%��]a|�-��<0�+ٞ���͗��N[��%���c�������H�b��-E�T.ސ����տ�E7L�]jX��e�w���r�Y������ߕ��Ff|�����L�8�����
90�Y-5�7��r}�v�������fǈ+��-����W��_jp @��6�F�$��/)�F� �΂��������9�Ʃ��y�b��~������<���Qf~~��2E��8):)))3G+@�-"�76&K���K�5�� �:;K��'��O�%/�9t�����-���nsC0j��C�b[�55�P�ehh+ p^����[��t~ׅf��q��ݗj��N=�	4s]�D�n�\�K�(/�����;��,{��a�V�`�`|��nPQ�]m�$+�x�! ��$��e/�aâO?��c�{޶뾱~a� ���~��L�x��Y[Êx�DF}�2D�-Tw�{�T�u����P%�AA2q����o��kPJ��Ң�~��5�MJ>555Tk�Ǹ���I�)L|L��z�rX���"����(�/.@����4�Y������|���A��jV��-E��/����P#�2A�C������
(w�p���e�/�L�@�`�F�T*f�p~#hĜ��[Am����������D$& �ec�$&&�s�`Q}���AhƊ��3l22466������V��z��o޿�YQ��bW�:�S�P�>1�����xsj�GHXbdɣ*IMMRss��|O`��ee��5�h���&����%�����7�#t2�{!��wxaW�ڶ�0�y�~�K��C�i2[�I4^ �*=����O��PjƜD8�~߆�XlNNN=++���߿9]]]�WU)6GЮ�m�h*���ޯ����;g5W���))�5���>[��:v�u	��8�z��^�+}�(*2Tf`f��D{N����5!�9k�ݽ��#�
; 	�M+g��t`�#�ױ���}��%s_k�;<��B1elb�ի9�MH1=�������j,}�" �nʈ�56~~�܇),�7A��b[��>��َ"w��rw���('m�\�?X*:ZJ�/Ť�d�Os���ȹ�fT��[~|�o��p3�l��J�dxh��h9$:c����tes3Y��P8'����v\����@#��j>���e�vl��[��6�5dEcf	�4����!=�V������n7����E�}���p�I��Y¸�]_«dA�4�����|��X��?Hnoo�00��#;�A�c�φE���δ����� �X96!+Ƚ<9顯��,m�-<T�Ɣ@��~|����#N4��?!!�"����A^�޾bA�M�+U������Ce����u�v1������YSa`aA/k�L]�v�D�Pi�Av���g�X�G����)D\c�5KΆ?�cdw�#�c���d�h�odQ\�,�|`��Yɯ�fYnrr+LŸ~oo��?@���f'ண;�r�6����Ą�d;�e
�-�<i�9fS�������ŋ���m^n�V�<���.�.ѳt6����au.Rϔ���>`c��ׯ����x��*�
�e3`ؕ�_�999�ʋ����"ggg�AD����%h�U����l�Pts�&��7�M��]�n$+��k�5�1Sm��fH��(���s�|�����!�	����`e�;0E��ex^�{?\L�ވQ�π��<�jG�~P�ٚ��J��>��c�r (x�I���Fڞmc�Å��8iy�闣ep�����q�o6&�**��-0DzC�����3����bd���$z��LMCù�G��`

�w�8���уԱޜ�f���ÿ����CM�r&��L_�� s��4�`��0}$D���&��0ꮠ�a�冄��l��::�Maiٙm@�&&��+ojjZ?-�7�Pb��T����Z[�H��o` ',܄�UUS\D�z����P���?5---��U�,s��@����Hh���2����rb	���N?��DBzΧ�rtR^(	�a�ڕ�`�`v�T��2�E��ʿbk���*�&?�D�ʑ�5��j�τ�~��1'k��_�v7�#峩�e:�1�
Ǘ>�Tt���8����N2�u�ؖ�� _�d̹B��Z]���u��r!׼�������{>G��冐6�ި*����t61�h�7�uv��eZ�5TK���ׁ�"����C�IJJ���3os��s=�1�0_k{�PNCBBÆ�'n
 ��p`PA��u�O/�)��H��u�%���rFGA����Gۏ�ޞ�������ո��s-Q+U�=>J��]�a)�/x�B�V��3ڇ�P����A�_w@����e�b�A�+H��Y�>8uz��(�0T�m�e�&2���v�D5�R�.�oj�{�D-H�:]T�ћۤ���h9��O�/�j�3�ȃ֭3�]��� ��?����`aiY�qe�c|!~���*n]hp�/z������G��]5h&��rNii��^���\:��4���$M�J��3�m���r��Ԕ�͛��8����Ն�f��#I���;���2	����������e�0_�����5�pi\[�}B��|������8'��T��O��ZW�"��_��CMO/�n� �����7��������X��������ҟ��������=�Z��V��Z�'�i����7j��/�j+ݝr�.�DQ	�`}U<��NQ���F'&�-,� �,k0���R��Yq�,���t�b�B�'�]�^�A�j@9CM\54H���������w��]��T����\_�������L�0��;$��u��� ���300���S�e���.s(�i�f@���c����j�S7��)���5���$�C����pvQ���j����A����{�f7ҵΙ	����ATn��ˀcaq�a�L�<7
��v�N�x�Q��n�ZZd������t#��tɋЮ��:�6]{k<�._f��U�y�t�z���(��&���ϳ���}�
��H��R�0J�W�>B+���	 "T�4�����Jh�XO&�u�����9�Vznuχ{���+,�[��^#kd
�0�o���R�Vʚ���RPC�'r*�l�#�V!�Q<r����4?���U����]��<\3B�����B�M�I���m�.�M]��Ћ�~��3<lZ��;
^iwVw*��1�B�11�<>�7�̺�Zć�����K�>��<<T�o�,���$�r�H��Q�u�+o�:��ws�>:�"F5��]� �� wX�����/W�ᐲ� �,T?��TO33�6��Q:��
x�Jx�X"�&��/�#�����|�`��<caa�/��7���ɩWG�H^���%���L��.%��>;��i�A��
�9rJ��i�<>�mML���.px˯����"�(�,�O�P)��x�b���T�x�^����Q�P����a��5����-�.*�ᎅ�[y�o�v�~[���y9,�gE��P�Qd&��m�θ�EƱ;zQ��ի'�\�\v���nR��u�H
��L������tɍ�+���%)ʶ���������+�l���3��8�Ke���`�����25Z�oo�:k�@��z��BҪe�ĕ[�eA��<y�T��?�c�qn!�,&*5N�T.-t��A�?�g����Q���76�5Ov����8]/�_2��%>=���*7);����O^Q����6&H�ְyg�iN���g��iF����{�}'lj�*��'	]��&F�.?������w����O�Vto+��C:�2������<�8xǞ�-�< Fi�_-�"�JA�s�=��_/-�ېsΪ���-=X�ʂ����M�wۻ�Z��O�5��� g���G��.Q��������kJ
2F�;��ǅHWamϓ-$x�>�
M!�~���S�I]��Ɗ�ڿ�����0�HRFtܴ�%3�P���	li��iy������gW���׃��ķ!%���ё�G6�ok�:z�>2>�ў�TY��<&�=�.ub��-�·�9�XT	����51�ƷlW�)O/�pqq9\ٝ^��ܡe�<��h��m��<d��s�	.��?���+<>7�����H��.%T�7�&W�f�`�� #b^vE1��s��I��G,�q�߈o��]�(*��(ʷ
y?vRn����XH�[�&�|� �ߦ�*�%��7�7��45�\�uo�_�R��ˏ,0k'}��\�&�O��8�N�y�g�����=6��n���*1m�^i��=ݹ
�ķ�)�h��R�X�|�Ynl���d�����L9�+��߅�bD[;�p7�RD=���
�
�#��_7Ej%��t�Ϝ[�*�Y�.߲��������e(���YT�@�H^��Jn�������{�'��'�Qq}��q�����^���l�������I�e�H������]Ģ�K�H����ǳ��t�F�����v'�,��ں���>��c>O�S{��-��d,f��33�W�4"����n�A*Q�\�T��������,�L�K;Eߘ��\"O�U��9VH|m!Ep,�#��,R
�y/%%�q��","����$�mC�`W𥄓A|/�vV|�c}��(B���ab�Gv���GEu�NR��d�U��џ�`���%��D���Z jx����7�JK�t![54�������fs��G�Ǉ�[3j)+�W�Et�o�9���}!(��m���B�bFӿ�e�x(r)�ӗ�o����Y��4id�0��/x G",TWU}MJB�����������mg^1��C	A��vW�]-6��Q�lH���<
��bXX"#S�iY��7x?)���ŀf�X��)"d�Q�=RԬ0}J,���/�?p'a�Z�ec��F ��=DB>��U�8~�����FuU��W��J��%��[���kM��E�	M���C�����!�%���T��2c'6c�db�QQA="0�˽�uzb?f���p�1$=���.;�:_��p0��|�.� ڶ4��E:w	ʆ���Y��i��aP����7q��{��f�rX�~�sf������� <b$��܄�]z /��g¬�}H���s��@�.bv���CR1��й+cYJZ*C�&-�9�W������芭����SK �Ax�ώ�t�����C��|��&�[V[6
Skc�nΉ�R�\#M͓�$\��H�����F�ϟ��8�k�y����o��+�2�#O�V�$˿�gI��1<��3j�C"�MT/ፏ�/# �h�6E�OS�a�?b�ѳ�������+���r����3%�����x����5���޹����p��D���� �!���{�O����nz��,p�BS���D�p�i��y�޹�#x��ɩ5<-xUrp�&���D{�ϯ b�=���P�48fJ����U񳆲���i���g����j��w0�wA2�v,��C���<��+!./�%��=��Dш��z�����O�X=�ax֥Ί��m5?�\IdP}������k���[d���L�V�=FH@UwE�����ݥ�q�t�1�v$�ჾ�\�\�9]�������=�����$B��g]��Ͼ������))O���F5�s.��˘��b�����2�� ����t.A$��Q&�7*y��S~^>2��#S��8|L�[�B�vI��)u��_֝�-6k�y_���ɉHwĩ@D	4Q2P���HX�,_���Y�J��Ie��85�Y�5��uYJ���?�3eLB���\���?:��/�X�0ǒ��,�������OJ��ڃP��S}���x������y���|��<Q|cYl��� ��+>>6VT�Ԇ�[�0J>�m����)Jʃ�l��ſ���߾0p�i�s��*1w�����#�J�}���ޘ��l��W#I��Ӻz���;��G U�!���14��@5���*���#��$�'@�4�)��w�G
g����qL�t_0)b"N�]LKtt��J>��m����-`Q�����%.7/v�������������U����Y��45)�:��u�M���Q��2�-e\���S!�[m��ެ/K$>0E~�'� �AoM��n[R�Y;E��C"ZGԤ�MI�]��Y�Q8����̌�*�i"�����n�ǈ��O#��:aU��0Nv^.S �X"�qnQ-nN�9@�� ����tZG9��t|��ww?k���k�ڼ�&7���ٰ��W����l<��L���EK��o�{y
��/Y����%{z�aR�l�'y���F^�RT����ս*|j@t��]�hu՟���q9�����D����*�E����-�Md���$�L�#��Dt|���/��ȳs~�����Jݦ����&_{W�g�#��
���ka��rځ@"�Ud֤����f/ܤ��?�����ˡo���Hm�7|�/��Е�W�@�l��� �O�#�+�5Kۙ�����"'���Z���	��H�gh�'�!�x�
�,,�N��*��llXY4�kWO&�;��D�?�x�%*f�o¼�60����)@G�J<�#�p�e��ʊ��>��e����w1c���׷��ZD�v���������,9��(P�R��tNx�ā�x�<)�^���Sb{���H̅e��Ϛ[����쑋��0<ú�SR�ҁ򕒗�t�,j�bȒ6���w�"k��=sj�r2^ҔYy��"�u?�'�
��e��N��#a�I�����U\�b��g�����%��}�HI~`}A���)	g$ݺ0�e�(�vd%���8����1�p�����{e���P^���ɩ���W��D��Bsw!-V��|�����K?+R�!���ѐ�%(E���m� ���v�;�?������d5a�q�W��j
�����i�\���,h���O��T�;;;А��AF���I��!��.��l���n�>�/�H�e��oF�9�!��m7�"�etg��nxl�F�#j��;�D*��7@A�P�ߜn�SzVUUA��gJ�N]:4�$ߔ�$)u�u���MI}���'&凿9�b�pM���Z�X�d��a|�\���Kڿ�_�3�;�KMe��UbEp����o�r5yƋ��w`�HHB��UWN^'�#��`�(�q���ٳ�}Ǖ�=����a{4E�Î8��ߪWL�`�6X��e���v��}��dL���Z�ZXZ�p >h\_�%;��yP쑏kn 6"��j��@���x��,cM{{^�V�6���[��G		��^��((F=�JRYHuWC�V<zS?�Q�k��N�?�v��ll�\܊u G1�ʪ�hNMU(�`��~׸n�_P�6Wm?M
�(P̄"~��]����rOU�^_Uv�>�H�a����h�y�$��`<���a Kⱶ���o6"�[L���<��/�bW@`t�󖜄�X����3�	P��1�޶u��,�13�t������I����]�H����WUX�G�K)CfO�2���ǋ���=m|,r�K����dAKx�ƥz�Ie---(��[F-Sȍ�QKU�M��Ą�����c$��mދ�)l�j�H#O�k"f��f�=��)%n���N%����`�c(�ݼh��'��=k4t��K#���{���(,���bh�S[X^�;!lm{諒>4��u�N�5_&eL���Fc��s�����}y�ܡ�y����+�c�/T�$Q=�m�~޽YQS����l�m'��3�g �J3�<|t��$�ȃL�7 T��e�ޚ��,�0fX^��JY��1�h�j�55�G�B�,�aA�^o�ΖY��a�t��\O���#7����� ��&�`xw���zz���yMy�P{����3���v�YJ�����P=�׌Y������~��}R���Ɔ�;췹�+��B���B7K�A�w�?~hD���VW�+N	pK=��~��]\Rd�2��_��z�u~�O��v?�,m�}A���~A/_[�ó���7f�ߝ=�ڂ��Qs�	޴�z�w�4��s)݀X&��E��B_fi��T&k4�/�W������*[O
��gp	�W��L�6�G�p�.N{����+|�q8,Io�d�V����g^��3�BU�Ã����[Fѕ 6r�u�T�P���>u�xp.�I�oʮ?H�!+/gO�gF�Ån�P�x�9R�;�C�7�jj�!��J�&^MRpo��$"q����u���/��z=��?haaf�
�)c!		
W咮	�%�:w �2�/�	����ҥ�)~Q�{ ����P]u�������t�:�gM�׿��`,�\���m��W�Dn�ѱ��խZ��$�(��H:bN��-e[9�e>>����������^Y �v����JK�d�<y�3��	�;8��o-�P���[j>�-��	D{���%�{�ja������k�f���rQJY D�D,�dR��p�h
?�ػ������o����8q��U�&�&�Ӝ��r<�g���~��n4�i���0Av�
[��p�Y$|����m
��q���4���DGGgMl���w�3����E-k�%����޺�����V>(���JlQ�K���B���A ��^[������$�l\ˬ�~���@�؊	Β_���G#@M��C�Gw6��n��#�j�k�G���3r�
h�V��0y!���?M�!����6���_&��@kJ6��^o����6������z+���w${���&*�/���\�^�fĆ\���M�;p٩��ģk�:�V��<�X���5�g�����%h��d��5Yq~q�31�q�ת�K���@�nJ?�J�UK��\�1?	�D}��W=�����ow?�����P��g��b���1�&��T�w��2~U�����a&@-F	)������K�tH�X�f�,*�#��f�m_c\g�o�|6ɦ�ֹ��o�u>L��FA���N�0]\���S���{��E4�//��r�Rm1��*g8<�{���4�Dgar��ܼ��J'�"�~{�v\����,�A�e��@�ϰ��/$$$�gO3ꀛ���a�S$�d�X�Q_��reb����c���#�J��W_����Vd�:)��%�b�ɮ�K3.��D��*�F�9��J|��u.ZT֐ >¨ ���}h�]�4%6 �~t\b��kϫ��6~��ݛ���aI��i�&�9�Ӗ*R�����=ʭ+����r�`�˾��ѕ5R�Yg��}鐝)�c�M
Q�K�j^Z���g��a��pglpU��(�~CeZG����ey����%���b�l��Z��z�o����P�e�KptL�R:ҁ�����O$:�2uƿ]+(:@�W���ǎ�%�l��g'x��d��R2���V�po�8�y�&d	�����(b�%+�'
&&bR�PKe�k ѭ��S`��2�;A酷����Eg��͍��_��)�kR��o��;��23'���2�]<Gޘؠ�M>Q�/ɛ�]��,��nBl13�~��;��)�%M �0J�W9��P},rCӿ&<��h��w��G�?�����S����NH�6�Dpڂ�J��Ą��l�������j� ��X�=`� �؊��s���&=��ߏ��q4����U=>qx�f�\���ZUI)h�^��)��X����߲��Ob�p�҉�t?�>í��/䴋�Q�F����m��T�v�K�kA����H����I%������~�?/D[�/[��uK�(*�j�wkj��H?d��+�9G2�$��*�j��d���*f������Y��?�c�	��H�%�!�1�������@?8�*�L����iX����V�H�$e�K#��7a*�k��-t�?[����>ZW_�s��\Qۄű)`[4�U�ٖ�9IHH����%�v4��f����ƾ���r\���>?b�'P���C���x*,���v�-hZ8�4���??Oz{{��m4,�O.k���U^��!�9�������'ӹ��3��m
��!���_�͈�&���&�U�q��
�*}0x3F$\(߻2�*������C�&4��=s�n�;��W�G������z�ɱ?M��߿�@��@�}��W�'�ϟq����
�����jNp�6{9|��=���R:��ۄM4b؜OF/2�_( w��-J�G���;���n^��R��QƮ�	(��S���u�����>-�����!jp�h����qgg������kb"�%������'���ss���K.�)SnN|w��<!19�o6�d��T�$��ٺ}V�)̯���#�E�΢yia.��'!]0I��`���k�}rėTW�V�j�h�����fb
���W�Ie��я�r����U8����h_�eJ�Q�[\QW��T��X_Tt��G��L���
����M�I0϶�vv����گ�"�� !h���r*`��#$�2"��(R5�P2��0�J-�W��o??��������_m�� �L��<��jg��r�̻��t#��c��)�QZ@���ب�	��mѼ8�p��I�A5��$��9?��I-SUyܮ����k�f���֔��3�ܫ�?K��D��d��p$4;��O��C��x�/''n�yehz�kS�Ǜ�1\,�aK��	����s����4RT��&f<�l>|-�{�v�3:j��������Aq>���F*��!mƣJb���J)��J���
�+�n�O<�Jv�ڟ���a��M��}�FɌ?�?�����=�&{IPVv�6��9�k�쪆�E����㶁/��x:K�) ~!!0(�9��a /���[Rb�>��"s#G��O-.�W91�?�I�K��};!Z�g���嵵U:RRRe�uww\?�`�di�/;~D����R�b�F�����\m����`����g��'�;��D+�j�"�@B����X�� �u��Ə�꫚��t������S���պ�}�O��l��'�Ai�0ŰF��k�'��F���,$����hTI*�ʞs�`2�1�Y��Vq�$s�� Z)�K��%�=ϓ��}�؝�@s;�lRG�����wq8:��gffA�1/%�_��%�7"��*��ɶ=�A�N��bb�f�ࠁ�������Fbp{b��V��+SwK��ӫ�@BDzIx7bb#kc���xl��Y�`�ݴe��*v�L�|$#�ڦ��*q�4�?��4���s�9>5G[��?��1:��m'��XM5��4jl[�m[&Fc�Vc۶͉�o�|��=k�ｯ��>g��s�I��|��e^(�a�w>�p�l����D{�`x�A6��ݻ�W#N&̔�?:���}�a-��qCi�;L~`�g�.?i��6�L���.��`X�:���3�L��hv�c3S�Z��a�
uq�v�q�d����q98�4#i#�s�)��;�L��_l�Z/Όpċt�\��]�J���Z��@-0�Dy�����t��c��ں��r�(�����C[�Vej��ɧ�<Ȇ�oφ�Ym79�1�Q�hG@}
�-$0{{��B�����$K\4�Ѫ�:/��r����H��~�yƏ&"�������D������Qn��Zس��F���-]:M��޵������ő0I����{�2�A�!�ZL,*t淞Q~t������WG�<NC�'�mQn�U;b������f �C�?!_M$� ]4��G�_�vuF �s��n�\X�(�i	�N0�n���כN���R&|�`wK�MSacۛ����y�,)��k�n�<��Z����{|y%V��@�@�u�p�D�r>��dN�����s��D���}�}������Aز33�\T���J�4�6��C�+a6(�VIVH\�![W��z�nȫi�X_OL����_����]�!(�K���Ufn�������@PUT&b�zz6�����S��Sd�tggg/ʓ9�so�Çs����������,�+�ֱ�W��ȅ�����/m�Y��ق�v�����\��G�\�����]�	�z��!J���;1c�HT6��s�?�'c��Vv^�\����=0'
�U�XYY���ZG�("�f7��̩��xнx�M�gb��U�ߝX���e�q��,O_s�y��� �F��E�h�(W`k��TMds�W�2��]y�D��������B oD���$��꼽����OJ4M,���NBwJ��ԲTB@���T��790>�O&�C���d�ʐ�B�sv���S�f�ߓS?45a�WS��˅�r��� �B~���yp��IU����dIm����"T��Ftu�^:\��ݲAC�9�QЬ�ӋdZ:+�4r��NJ��(�{>{Jz/�344${��ʪ3E�X���s�حY�K�	�]$�e�:Ȃη�Q�6(R����q���ޮ�{�/�G�'����٥��z2���	�"!\+���~��<�OjU�	<ۢ�	v���z��d�P��o�;�Y�,l�٣��X�.�n�ŻxA�����_N��
F w%����
���D�iϸ	Bf����e��o6{�&�{s��p��=?�c�rm����*H��<�+Ec<��":��-D}&ʐ���3j�t���z=)��fow�3ֱ�!�����=�Ӆ���X]�w%U��C
ŗ�m譼���S\C�At�����;\˵n�8�ک.��]YYf�/J�f�H~y[��䨫Z�ۚ����N�0��m�}��g�CRX7�~�|���/F�ա�@�c`L�U�$e���l\?,,�^z'3�ax��֨��Z��K �_�Kf&
ER�G�:���%�k$��o�pgߞ� Q�Z�3�̑�[oN7��uY�O���K�?g
ycSa�6`<:iW�Pa �; �p�V���`�z�J���~�ͯC#T��S�����'��İ��'$dp��<�^�QǱQ(̭��n�lՑ<j���BX�Z�Dq�;����f�T3A5�Z����s�Ph</]���|�g�
Q8e����g��P_�5�|`?��BMMMYU4dZM�H>&�3QI�%����x�9���Sj�NZ�ޚ|����16�&�i����"�%���#�5J���1���],y�<�"8=��5�_������YX�����5��H���'-ɋD��*�L���@x���(@g�b$9ia�@a]W��;u��6���X���L����<K��\C��{��W�(��b��9��Í}���_$�u��gRR�ah�p���㙌* ���54<e�D�7վn+���Љ��`�^�\���'��H�W��ܱ���sV ��振/��/�32>/��(�j3>��Uλ�����ٸ�{�G��N�9��<ϭS_��E5�����+,�g�@��;BC7�0�u�n(�P��q�2^VP�L�I�n�7�Ppq��,R>�GQ;ՖMvU�V�u���Ҧ�E����Z3fr\B�E��G���?m$����|�ȧ��%�;o�:B,�M�F ��y�H��Ƕ���$�c~�}�ob���85JV�#��Ѫ��As�i�$Y�f��V���VP0[�8|��Z��d@c+{�0�'%OL3�+&�����TM����N��'sj��w�9VN+�S�đӢe+���R�-01�Tܒ��������1�O�::��5�{$��*.�dK���@B�4���W�$?���I�5�!h�vy�l��ep#�J���#28�<a�W�P�SI^e����%�-~�E�z���� ��>xbt��5$��'�\�����:C!��̬�f�>)p�\�۴���`�p�g �묟_`e�.@TC����8.IzK��Ar*Fw��/M�����5֗�p�{�V�)��	�񛽛�Jd�6�N�pS�6��qr6;�-A;���7�3�ؠ�����N���a���ھ��.M�$��L��S�I����5ګ[���lL�֭�*%DPK�G�+4��s����zr�D����������V�d�U*�4G�A��̡���N�����I�O�NH~�ޓ%/)կ9z��&�Uh��ucpx4ҖU�6�6�}�SGTY�koP	{<5�ݰw1R�0�N���'QkԕϐWѩR����E8�k�t��\�6��+=y.tƕ�.�����*�+��0���� ŨU�3sX�+ʞ�Gbq{�=�t��oM��
� 5���Ɋ��r��5Y~YYK�Gm��F_k��}�5�?��t>����b}��1�مC���|,��E�9�gq���[[:ޔ�Eo����h�M�
;{�DA0���2MP�H4�a�j�LTH�U���i�h4^���P7Z.*��ݽ���Ͱ!����19k
�Y� f��_,GѦۿ�dk@��h�%�v�\HR���t�7鉼�T1��'� �aT�90�в|��['�9��Wt�<:J���T�Sg�K#Y:����s!_D�w6�!���K�0�A�1�TgZ�f��B"��������O�����ھ}�FJU)ַpp�]����k��0�<�1����\n���Ohi��;8P�%O��U*�Z?3G�����b[��X�RK\�s930D�e��Q׷�&P_���rF|�8��U�9��x6��C�2#���b#}�B}�0�Y1x�W��By��`���ajeE[��PR�jk ��/� � � ����$���H����
��L��t
bZ�� -`@Wq�J�>�.�*Y(� �#Q[w-.QƑ�Ig�=�$�69%�{ҏu��h���i{x�I�?d>̻����Y�=���a���SU�d�����4����[xK���`�MUɜ8ǧ0���ˮ�pm�Ғzy]�4]���`�gޣ����'3[J4�ôELv��K����h�g,�3���.�۳"^�����@a�o-	��q�ٹ����p�9�X�5V�_�n�����פ�t������Ɇ���**�$'|� e�%c�q��*��
5#�B�w[{K������SY~�Lhؙ�~=��-��$q۵x%�{d�(�k��֚e������ V�N��G{A�[��D�Fm��Z����^��@qk c���C�X��cT�e9x����(��6v�.epT��tq����`/$���a����Y�xݳ��ԣ��7E3@[��Y��ү&F�{�O�V�F(G�j����Ԙe_���^��8y�������[Ⱶ@���8���.���;A�s!��S�Hy����,��K{��>�%N�{����w���0�[��%Qʯ�V�f*4ɣq�]xv��Z���dZ��&eRy�3f����U�,�5+�cO���M�m�g�Y�a\�<~03{m~~ �Ë<~8&]x��H�L�����K*?_ka�uyS�M�nO�W�Ց4��l�
Xm�램h���/)T��e6��?���X��S`ϜZ����^���dh0?��O�Ţ�cO~Hy7"����5��׏9v���lש$I)����FO��C�4���x���IJnU�N��J'�1	��N����̘�8����S���\�n����FsXe����5��5َ���f��[<ǢR�eX��.�J<}����%�F=n+dXF&&ϯ�2P�:�q�6�@d)��e�l�j����N�H�NCu��HI���
��qs�>��IG�H�Ȯ�9�ģ"���)�f�[��Mb�!S��n�l|].�"f)ĊI�27?'��;�����݊��ӽ��|O!7f����@)2�nz�Z��vI�����`[fA��^s�^�;чM�$��t~`W���#�6�*������ִie���`1�,O:!4��#5Q�����1N: P�,��R6�e(9�=�+YV�8c�]|�b��+w��rz����&�)����&6.Ԏ.l`F[�Oާ��� ៴��)�:�	L�u�/	������C%p?#�9��{�Н8� |��`s �a=w�a�û����^;�/��*N��:�hn;N<]�����G���{Du��"9q�w���n�S�����IO_,�����<�A�bn����k�8>���â�;��Fg���a��x�2��d����Q��٩�f�!8Z�1?m��܏�A����U;�;Sq\i�j���D%���Z~m�s�0�A�ʫ$\d�
g�n
�{>5�@�d�dAWr +�l����5#��v����x�cGιKiD[�+F!��S##�$��|o�T�%�%1���B9�GcZ���ޙ��\���=�C���<�n�=φB��~��1�~��'o6eD�扙�b���~�m�I�j`��@&���ҳ�ǅ�>���+���
�'����O��!'��f�ʐ�fV���Y��'����t�	�:���)����8��|��u�\����è�`&,��[�����ܐxx��� ����TL��ɑ��A:8�O�KHRj��bg���5��p.�zF�������/	ӄ_ppTk�l�M-�������j	"�R�q��H�f?�8�z�-N�E�*'uӥ�y�:���w uL��9��wH�H'>��2�^gJ��!��Ohq���P�^�ӓ���3ϳ�%�+�XHߓ�h't\�q}�ڕ�B�>)��$ڷ�z"x�n^� Ҁ��5�8�^���n���T�\�H	Ix���´����{b'I��82"��y.�y԰��!��|��Uɫ^QcMB�U5 �#�;d-3��n���A2�)GB�J�-���V�)�8GA��Y���;�^���oa�G\�A��
F9���bw��H"�%��`�Wqi�b~H<nC_УH�vLM����H ��K�>{2���@�k2L��w`�xˈ��^B�����T_�SGq$k��f_Kz�4�dh ��cƅOp��w�[T���7��'^����2֣Y	���9[3�Q��g&��Bew�@z�n��9��:��>���љ��T)O*+�7�q�0AHA��u�~���Xr��M��3:��q�8����s0�l�)�DL���.��* n�Q8��&	��Y�9��<�׳�s�悖Bs� �1v��i�>�t�u�Ԗ��V��r�N`ƀ~;Fc?�}�j�>#������B1M�+����{\Z-�*�N��#��q�\��X��"��<R���%kkk�,�<Q��Ш9��y:"�1))_Q�c9|||�U@XX�&��-�2��֪tU��X��"{C2�S#M�hlZF_�sD0l��r��)�%�Z���)�`'gbZm)��S3k����Vo"��d<������7���y\�⚋�Y�`�:�㎁�sr�UeK~(���TY�^��v=s�/��_��/�0�B�gv�Uy��p�7���}Nc{A��XR�?������ݹ���w�R��������!L��M����͍�Q_�x451�51 ?���u����r�=^L*�wԧ�1����_bmo���'���Z�y���Kn����������~��[kH豉�'%�~u�6m����8��v�N�s���.Ķբ�����'��<3�q��?:n|���'E���'}�S�y�m�u݆�
7|�r�|ZD�ȅ�&6�eYE�(�,k��
K3���JP|������.N2���;7�-`�#�v��M��,�TΓ��)u�dɊ=z�'1�u|zh.珙����x2��KD��.���M �h4_�T(׀9[9uZ�A��v�8I:"�rS)_T��Îq�ޮ.��ƾ��y$٪4�MZ�K
�&2du�sN����[��'t}�u��d }3��Q}5m� _{�!�]�Z����_��3+�2mb�8�$���و����4����jE��ſ���8'���z�p{.�`c��Ol b�����.��s��_5��N/O--�5���*/�$]��+2�r
�@��!�!~
Q]��Va�ġ?,����,ܤx�嶥�<�ޔ�RB6^�s�o�?x �1o��e}n���FS��'�	ک�+�h�~�ҬD�F� h�qj�2tim��aԒ�ԐS��F1MMm]<FC�^{j,Q�B��,xӔ M�-$�!@��Rc?؝�pO����_�.��ջ�GfVk�]�xM.b�L�Fu �XVb;[��1��~A���1f��Gf[���胫`�<���]����u�}��������O��.~�����v;�ӭUy���B����[���y�,�B���p��ʩ��fT�6����zuW}���ډ��xEa��0a(?6\d�S-�*�8J�n�2�I_���̎��O�vo�2��0�<4�q����M2||^����L+�0���i�uR^"�:���Yﶯ��I�^$I���]R��m�?�@oU�$6;�)(t�9�zn�F)�ڲR��~nk�E�%l���$�D�7Ե��H�OQ����ؖ�;[�h������H��z,�%ئ����͖��r�L�ܧ�_r�����=�B-�/"?�	ñ`s��u,��,�A
2l����#N�k4��(�B�`�*�,̸��V�<M��9ޟ��d'���%�8�T�,ϐg��@vY��Äq�m�ɂ �V��ȇͬ�����sٍsE�Œ+1%��v
�c�S�a�i���޺>L;�B�K�ydHS���g �݂Y� %8�OQ,��H�Y�5�W��n�viq���@�),*�Z}[�]�������'�?�)�J��vD�-m]b�Kt�:�v���[В(
v��R�����[�|�*��u�`�����M�q
�>�it�g�?�qE�%�	E�V��]<l���u30F��+�+�Ļ>�� `*���mr�c#M��H�#�E�=���?u��K��d�/��i;��?�ڀt�Z��/
��^(�FJĞ~�����e'{�rs����� h���Y���B�H1�����oDB���%< D�gR ����#��H���k��# L*QXO	�/7B�Q�[>mI��V��Nm�.h��I]����1�����Fa�-��<^��Lw�o�h��~�[N�d:"=$6�/��>��L�L��a�5%t���4�b��=��cL��a��h�ǎ �ιSm��iPOI����F�/�ZUN���t{��65�ޟ�fT�e�:�_8��` 0��K�0R �ī�>C������,?QRURO̤�@�<p��㓽�Bu�+���ޠI>����m��m�'��n��Z�f4](�����Q�yi� �5�٧m����Rp�OhaP&HV��u��H�#a�t:c���ߍ��hD8D��ұL����y��o�&a�F�o������p�E ��ɓ.�������;��2$���'N���b�@��w�|�G�ӪM(��[���mg"d�����S��#G���EL^���������D�� ��`��N���=��e�|�2� �Z�
�})��8%����&�ȲmO���+��@3�	��A�#cn�=����m{[�"U�A�Zn6��qh���R�<t!Ht[\z���s<�mc|nIn��rS�㥵c���8������LP���U�4�A��g�k�)���O�TI���h�a�i�3�[��ua���� ��0PH�]V	�`��-���]�Ku�U�|���mU��X�ཧ����dW�߈�ہm�C�l �8~��n�}}kֿ;<`��^u.¤hcu����F��fB�������l܏H0�t�Ծ�bI�Mvkv��Pv��]�+H �d��۴�LP������7T��;v�D1�+�����A���<5;�$g}�����T���D!(P�x�Y���)Ȳ2�M���*���#�����9¼�_oxe��19�k/2���3��G�M�jՐ�-�iw���?)�>��dz��0-<����
��NdȞ^�x���7,�V2�CR������ھ��qv0��|�h�";��'H��ʐ:��Cm�ϐ&x@�j��1�-��{K� �7@��o6�	X�(cּE��<|�dP�� �7�@$�	�����>s�n;�كZ��!Ϳֶ#jp�>��a���3�RuXk���%zH؋�]��qI�#�X�o��6�V����V�I�GQ�f�I�ax��e��d�f�L6��ZK���P�/ P�tC�R`���o��ʂ\r3h���Ԙ����:
4	8m��`ʒ"ܛ��LBLY�8��|�1���~�y{��B���j;х̊?�,u
�(4gTH��U�n˨�U���.���GY�� y��S/����N��F��(�}��٦�� �a�f����8�y)2�j�0a͹�%�76�`�ȳ��2r#L�$�=3��n�;"
��L��a���)���$A:a���)$�ey�A�	�%�ګ�~cQ��kPe��UXL��G�*��&Ͷ��iEْ缠�0m72u¯ə,�� �~�m�����ŞYP4'{1�7�Kݱ�`���Yw����"�Rlu�KK���'}���>��Zuj�&U�� eжՈ�)h�?�F����i�*�С%���np�;��aΚ�@����/"*L~�a4?���T�9�����N��N+Z������v�s��8X7���+����v�W��nK"A}v$�2���)�hg��4D{�V�N���pJ �U�$ �І���4��Q���ȌVe�V��h;=�.����GކG�M7ίO2����m�s��#�uI�6�#�߄;�]\��Y���B\���q�h��}ә��S����_?T��N�{���������P��\�tj�0���蓺�c_u��P0�3lӼ�s��s�g���oƕ�m�T˱�d%C�C�q��庳�%*#Y�Ln�w	���$)V�Q�f���n������w�_�����[pE��l��]��T=��?�w�R��:q�w��k�MB��Ŭ+T��.�bG�o}�v�<q�};������F
�R)����#���g��&F~���v�]ik�X�0��3���<�ɰ�w9�R�ݚ�P��	���0#�6dY��{��L�?�$��L? F�`���Ռc��z#��b�7�'SQ絉+IɄMo@�67�X��a��nt!.���ӏ]Ѣь��J=ފ��灐VB�ؤ���nO����OtI��ࡃ=e��
��S-�V�I$�����L@�7i�,o<����ࣧ.�?j��̡|����������K@�D�<T�JyfQ�K �
�&�j
�2��ח����>��@bWT�*�v�b����c�ۤ��³��&Fn��X�����\b��Z�>��Sl�Uڍv+n�? W�m�� [{{�ti������ 0��7� ڣ T����wi�B%�ѝ�v��M�d��W �E�j��g8g�iG�K�Gt�/^���$!a,����6�w�f(���@3��:o!֙�Q_Q��Ѹi�vg�Z�oP�WB?�Wr~�d��L����:��xZ�؈d[fOcrSX͈sv��d���?��3`߀��FªX��	q�>�7�%�u�F߀�B��y֓_�\|bY��{L�ba�5<�V��Jy���A����j0Z���� �\W�������,?��iX�7u��ʥ٣1[!-�܅�ԁ$����LQ��$���Bug8^bn#�y{[Y�-�7B���B��	1������	4}n��CJ7��K�z��rhƃ6|��
Fs0>4.	������ގeÖO�d�l�{�����h�r���
�h�m�����;�s�Ҹxx�h�vv�s��ژq~G�?���>��H�X>F#C�����	��d��F��=���.�Q_��-O5nB���V��/Z���MLz��ⶦ�H>³�Z��F�KPpp������dDʔ`tH�|�p����E��_��Z[%���%�	�V������_`c˲M>��`�g��ej������L?{��J�t,J����ä#�H`ŕ��5Z1�mf��,P���h�G_���������e�8ol��!�>�֫��
�~
�7�qH�����s\'3�ke�k���ַ�����Ѱ���|uP�1(4p�D#>��G8u��_��u@K0{�xܶ�cq�5QMF��&i0N|"�ڞ��,i雵�7���E�Y���{.2�F�����,��u.�����ێ��(�v�|�հY\lW�o��#H��l}�sf�ALM_�M���ꭥ��fbb��1?�b/o��t�m�@��M�@�����䬔���_W����L
��%�I�JR*�W� �F5B��A�W|�}��w��`r���+}��8�wW��vb��|��%a����b��Hñ͊ԇ��s�ݟ����'R�.w?��_�Hp��39�ֿ:ӑ�H�����8(���?�H�N�I�W�5~�%�g�������"	��U�?��!9ϑ���x+��ȔW.|g�M�o���G����+�hD �"}�gR�iB�~�ﱐ?�Y�jrr�]�R��I��5#���墍��|I�����������"�X��,���x[̦��v`��;p��Kr���.��bP�>���H;�cs�����X�q�j\�� �дZ�l�ڂ+��I��+T���놢
�[����X2h(���7�R��q�Y����\�q;dL���]�R���_}�{:�w��E���)̭�O��W��y���s�^��y�� gZ�OD���cc[X��;t���U�P������՚����;��:Y�0  ���
.���6�d���/9��A?�?G<1N@x�\��`9����cؠ麜�G�Pn"xvG>{+м��G�`��۸��Az��:/�K�u���|}�2�|���{�S��������1+i���Ĭp������������ �ӱǝ\�8�0y���5���v���FƊ��}Gr�D�]7.{�X79�}�fy~��$�������2�SKH'h� D���H�\��f��m��i^��X ����~G�>���=S��Q_�J������	;��oٮGYU�N���H\���B�Mu�U�|1�����_����S�gK���K1��<�P<{����+������)�3,�M�f��u�N��L���e�ɦW��T�152�a��H��x������tf�����R�2Ĳy�Dp�9�Ο�G�; 3���b2A�do?�9¥���˰?nyt%6�fIZ��[�-��fȾ�&��3E:�>蘡"�#�D�I3�>Ì�{�;���@+G~~cG$�ȒY��qv�&�!�у5-VvC��7C��2��*XW03c/	L����ٵ��t��cN<�*��w3ꌌƴ�:�!�7P$z ���E
�����$?<�����::��2T�3ĩ��ID�`h���Ѷ��U������H]���R<jk��7��[c�
�w�ھz*e0��+a�)�**���8����4�����\�� �-�:5`�'?�o�\N»�Q����p��Ķ����ʨ'1�D��0s&� U��n���%A�����~$U���Ns�._�6:z��}3�h�cc\~��K
Ĉ?P�n���W�Ld^U�����O������Gy�M>1g=�m����{���tW}%쥭����>1�'eɱf3��Ֆ{oQ?��	E��>��7��cv��ۚS��~�v�2 A�dm0Ž����^�e�C���^\Z�vYU_f��&����x��0vf���x�Z����y�͐�ӺGT+&6���F��̟t�>��K~�'3i>j~������&��<`���\ט�<{�ՙdy�)�����p�� ���X�Qha�5L�'��
���ߤ���_7�CmL�� 0Ily���9�7-/�x)O���?}�8�_���Y��p����#��{��-�W�C��p{��b�yC�0�^ W_(׆�������B�B���AW�W�Ŕ�1�S�`�$B�Р�=p��!�Aa��#�t2��i}gǠjRCL������-)vt�斃�H�5ڔȲ�ߪ'�?;�t�&5�G�s�67�?�_K������a�x�=��9�$����M�f����m�m��a�d���I�ıw�t�ǅ��B�	
��d"���Dk|��z��t�W;�w7O��1�4LQ#|���<��u~�q.҂��Zb�d�;w�%�)�:B4�-��c,�U���,�X�{<��N�����Y�o?%�=��e,=����$�Μ:_��9"�i�&��d �0��TONJ�=dN��u3u��@��c��3=xh�{�����6���|�@�B�OƸ(�8$w����<�	�Ц�̬?aS�τc8Y��v�����J4���R2|�``�y>�R���U������6���=�Z����\Ί�0�7�����<ɉ������Yo�R�.5fz��V$�d)^n���ْ82�_�;^��a�3���!j5;m�~W�D�Y����e%��?S���U�>l������҅(�>���U�ZY�L�\��\�˸���T�;�����1�{SG����?���Gh4L��$[�-)P4���F�⌜�`�0��0��y )2��eǻ!$����i�ig7������C��f�Uˎ�L��<�L����3a-��I�g��3g��+έ~�皧[7����n����W ��_�܌�y�樊�����U{��w@.����UCC#�r��_eNF4��ϑ�᮫2��4,B�~e��ˎ�k�;@wOdD�-�3EQO$�c��'CrX���#�;m, �inI�
�uN�i�� �s�vN��Ĺݪ��T�� �1��� l+��gߕ*�ː��-5 1���|c�����C����yX�)9:}����^��S|\�~��й�h�`�����߱|"���9�����9K8��p��\����S^��k�[�w %V�3w�Y�H֚�C��8�����!��A2r�f�O�%�#����ֱ�Z���4`Aр���4�V�e�I��**��X�C`;�/jCո`�;��15I��鵌��ӊ��:��\��@�li�	l�:��Ｆ��FF]�/u�]�"Y�y`1~��Q��N�sAL暃:������z4An�J&(:u����;/Ք�$y��N+o�1tE�Iτݕ�������Q��F?X�M��Cl�y����_-w,��p�L-��b��O0f��{>'7[L�y#�A$������1��@cQ�n�U�^$�]0�I�K���\���!e����
2�!+15��uǹ�k�M���>.Q�D�����	����By�����+���)	��ri��?���#V���Z��{5j�M�@Q��A�,��y�f��@�6��:���fĽn�WN�	���f_m�J��w��p�}�'..b[i�0K���t�j��^�*`S�%�<��4�w�qq����;y>�zx~��}j��M�@qA~�C�|�d��JBo�����	�ZL	�H�7�݀��;C��6��|��5�9����T3`������9�X�¤S���ơ��iXX�W�뉲�a�%��B��f�.3EDF�\���ٲ4�O�>��B�I�/�"�hRڛ�
���lmaI��"��ѭ�y�嵔]��@1 g���zq�5�c�Y��$�4���E�xF��q�/r��r�f���_��6��Y��ڝ&��¿�^;��k<~M<��~~����L��*z�,����~��nz=^������o<�]|(6�Ъ/ZTB(�#|Z�?��wK�����8���f89��z��[&dJ�=-L<>�H�p���a� ��x�F�{���+��\���s���#���M��}�-�䲐
f/�,e���Iz	~_(g/}�O}f?`�9�L���X�G=abb�%�X0� ȣ�M���ss�_�O'R�uV+��p���l�/�$�b�\�f,K ��h�]�~2�]=E�d_�ʣK���Q��R�ZPI0�rL�7�m7[̧s%�P}��-�"0+�==e&���5��m7��Q_v��&3�6��[mq�Cz�:��2U�����\� ���(ק��p���Z�<�у1�ެw;��k�:q�E�ϓa���˞<�	��&�ɽj��g4�uǅtN��Bv� ��\����#���2����妷�A�Oт1ƿ�Yn�K��hF�Z�G���ԍ����k{}{��_���{O��KI���æ$���V��ĥ��}.��/�	h,E����u���gS��Ƴ�{���o���<�����3����b���� �?URX�Ϣ�(�a�W#���D�P=!~Q"�����'6�,�؎�*�RN?{|	����������@�q�	l;���y�;����ف�_l�����-?��x�qv5���XK����(x_��ߧfдBf�{(N�C�c�| ��� >~��z,���8��q&�g:FG"C&�Ÿ}��!��OF�
U��A4f�7��)���cO��i�o������8Y��sW�-�H�����Z.���5m���sK����u��u�(���9b��J��ʅ�`|��_��~�
��TzԨ��iԦ�ᡠ����m5���[�V�:8����;h��S�߆N�ڌx��u���)˼�ֹ��I�����E
r�MP ���ն����9��5����)k�>nU{���ߦ!�)8�g����;jο�q�%�,���K�*�� |V�V�{�zW�4�G�E�p�F\�HI��������E�W\ͫ�֢k��% ���C�mO���,a(`�eV���c�0�dDD����Q0�Wm�R8}^O���`��vi�B�0$�N-.��/Mdɾf��k�/0�Q����=���a�w-��p�%���x���_dV�.}iS�.&�""#E||�J˪�_Y�r�lQ�)]x9r�{Y���/�Y@�>(xFh�Tܢ&�^9}z�,X����w�>��i�k��_Ic��>�7(�V\W|Ѡj�29��:?p"�X�y�hz��O����O�<ɾu���|#�'Yۤ�P��/$➆1���B���|����G%�E\��.=vkjB��\�x��bߤ_~g�޲�5��J��&G��u����.@���@)OUƹ���EL�Ar��qb���Y��6
G�02��aL�9HD����񁪾��e��W�
J^��SAl�
����觜�9����ӗ�B����OO����O?&���\�A���f��a-�h��S(=2�U�/-�j�-���å!1�cq�18g���P!&Z�Ƞ�=��x��Xse���{�.�wJ}�1���5 �k^{t��y��L�ͽˎ+�[GI3ƙ�g�X�~��:)�v���S(+�(���O�_�1��]� 8˳'	2Qx\Z���E��A��7YYj��F�� �ڶ��<�g�goNw�����?�x��WX��-�ΙPּm�P ��m�>z�>ګW��5t �o�o(�9��5��0���$�R6t5�~A�=��xv�a7=	�_�k�P�fY�ܜ��^�O����l:��K���Vs�E�{��J�����S�D����� %4D��ATW3T����3dҤ' kS�����0g\��.[�5r���Ǻ8��o*&*r�]��>7��M�7\���Y
EE�ؿ�mKM��θ��2�
�����yHSx�����h�S�e�b'��8:�i�mn���g��z�f��n�4n�n&�Ex_���[Q��laY#	�o������.]�����05 M�}�Қ5>|t�xw�?ڽ��JIn�F;v��������&��z[I��d2������q��x�=�|��D��u�h8p��qI)򳳆���[��n]��ݵhq+�^��Ew�x�+��Cq��nA����;����{���d޽�^23ɬ�[T�4:mbeR�%���W|��+|�v7/W*��Ʌ^�t{\s�EM ��ʵ�_e����1U!��qW��3���u�ƛ��<��� J^��Vc�ި|]#'�^��y��0��5<��߀BL�ٸ�uBh�z�D�����U�h��R�K�z!�G�h����O��j��
J�UX���ni���]Y���F�Ek	;�o��1�d�	ly���|��E�EV<�k��E��ed%^n�H=�M䅵����?��y,-s�^hq ����g�tLw��nj�ډY�W�Z�GC%5C�	a�I����v��[��#�}�k�t�}�I<�V���H��<B����q,�S�q�H~Y's$���ؚ$�<\#C�]L�� P.B�/ ���9����J���jF��S�Y<*�b��qc��9tɳ��gCڈ02њ���M������k1E�':���6]�^��k��Dj�8,�����kV����?��͋������Pɗ�N����ñ#�b�o����wX�[08��f��3�s�3��3h(,�g��Co���/���G�|������\r���TT]������A��q�@y*�L����w�t�X.Xp�'"O^Bm�x��l���_[��;����h�J7�k�h�{���A��b� �uG��T-�g����2����ԫ�J�U������5|�;��C�I�h��Z�|����#��F�h��m�F�<�Z"��
�����vՆ�$�{�g?�<�ab��Xu�,,7:@⫻!���T�Q���a�Q��$�m�J�^I�����JM���v�Q:姆�,����Zg��I��3ʔ5��MID�E	k�{P�M�(��]���윝�S����rÁ�w��7u����Z��L��0t������SVH�$i���OS�y����XP�𮼬���e�z�Eìx��=Nzc�(�=֌�9�&�b%ʹ�j�.4UY��Mo������ݐ���5�㑩{����CqA]K����ʡ�l� ��4	1C����I����rj
�$�Nl�z��qG���|_�����̕�R�`^�^�%4��@����!���M2{�l٫��z��2#�l��\z��O�$.3rf ½�ο�顺c�d֜�ΪF��PZx�J�f��GGdN�-,��[K��łD�m2�J�m���-{�0���A��`>�qמ�e�Y©���-7i/�=luG!�Ց�e�$�%�U�����o'�V,;�U=��	����������$�,��]4��_N�}͘���hxS( ���?���3��"0�6H�Q�u��+/�~�7d�E¬�\�GQ�����"�5vb�%�Y�����i�7A���ն�8���۠o���,Ϝ����M�|.)�m�s� ��+��%�l���-�w�o*�I�{�B�ˑ�{���<���9�C>�p�?_asRV�rpً���A"�@��
"Q�rD M0��z�v���-�FtW�p��^��bl��Nm4E�y�{���J�`~|k�N$aa���$���Go��� ���AG<��
�����x�Gx����`�W�G����LS�=���+e�Q}��^5.��RI2��?��3�Kq(f�2�L�4<:��ۼd!-��1��x�3d��m���	�P�W��tR��o����/S����-����65�ǇN��S$Ui�Q�G�Xf1TYY�KhK������B����eZL7G󛗏�	���8��T�W�o/ŝj�Wrz\��c���ك�x����b��e(��b#,��]VQo���v6���}%��Pyk��e�X7&l�d����϶��0쳷�����1�0S�<_��n"1\]�ׇ����vV��!Am[pF��Ö)	A {�0�%��U�f��ۊt
<µ��r�V�Q)ݽ�bK0ccP���tr�ӛ��Ҟ��g�2����|�"������&7�a�"2�p�@��;;=�����Q���bc�ˊ��-���� ̟�bCpj8��e�a��P[�N[ol��k,mQ�&<�1��L��cPeퟐv���gg�U,� �/Fͮ.���e>|B�	�i��
d~!0��k9;�˲����C��2͢���T���Y4FyF.�m�u=o����(r��6�RA�m�\�_E^�@Z�
46+�����0�fFY"*�^�3.+���L���˨�a&�*?�\��t4�;ȗ�%P�����<~߷|2���ȡT�&$'�6�7��mpa�	�+���i@�Ryn��O�]�)%/\��}7b�6a�XĢ��_��;_v�V�޾�3:91�fڇ
�]]B�hE��ٕ��p��Ř=�]\o��q;���<�-�O���>�)�<Z�V�d5Nk��o�m��>?}�7�IF��8���K�̽�nA��Ջ%���P7'	�>�o�\G{�l�d��m���z���(H�ף�]FOݛ�L!虫F�_�(��ym�l%
@�D`��@f�?</�#�G䚔WeKZE�����Y���+b�@�SJ�Q*8K� Y����즅ǭ�߱����n��f^�Һ$�� m.����8!g��*y���nOVMfC	��jK_�:��ţ�)�L㦖N�CC������s\�
S{e�@;���E�P5��i:�v�CU����B���m`��{�J�9M{e��Z��?/H���|��J&����.S\�@��ﰴ��h)��ι���ء-�ΰ��u�z�u�f��c$�c|�h�ty*����=M�y��H�8k�7B�0G:M�E�7�dB�'�`���P6]�~z�`��׏�������]�0�������0?u�]l�R�V����&��,8{A�J�ӕqt�Z�ٶ'l`���d���?��K�l�Hzy!�%�l���G��Pt$j�L����x릔Q�-_�8��l�g�W���/!�A��Ʒ�;ݜwa��gR�2+"���!���|y�(j�o/r����t���I �hu]�:t\�C�-�ā��G�B�n�)V�\�\�?;+�*�n����ILx��#���LN-�/I���N����q˫�чm����0�*�K���~Qw�����޾m���ia&�6W^W��`����Z�������R�Al��|��a���*j�%���άOA�c�����t�y{� =�O�qC��z����e�562��fD��X3�t��U��mT��I^��O~E A�&fq��~~��24���kdȊ4h��C�uբ�9�������$5&΄�~�3��~����-C��/����n�W���ףc�}9c/�<Z���2�?VO#���������6�h�}�S3tr�5����e{۹J��n�q� ֢tX�l�m���uU��r��vo�fp���}QMe������_@f���+�'S��6��K?U̝��Τ�(���P;���\no�j|K_S���	�&���ߵW(���!'q���vj���-s�wuYe[ճ��I<����>��Ϯ�{�	JT��D ��<q�����:L�������KX�/���ӨK�ˈG[X���IXZ�_܏�|���aQ_`9�5��_�W��������i��>�n)����&�!��Y�/���	���U8sx���ˣ�K\�9yv���S:��|����|����\�9����r�f��L�I����:^.���#�I�K�j�ʰL+�A��w]��o���ۏp��`���-o_&=O�)H����8���و"&2q�X�j	��6�cN�6�Ľ�����	���f|ʤ�_�]`���y�����:��05�8Ofd}�UG���ҩq��47�oƯ�;W����8@���l�RX6�?�q�K:��Q�a}�� ŵE���T^�/��G�1�;�%KR�^�!�\�`-�ߪm�=�m�g/Oi_W'/��C�N}C� Yr��H'ahF���(��u֪s�=��M��3�{kjjZ�-3����fjM�����y'Β(�����g�@^^Y��OR��1�ֹ&nq����g-���|��|��2�[O�)�٦q��a�4�B�HRao��c���LG߾�q=��tە�8���
�f���1L��+7 ��r~ =5�[��(<0�o_e:A����ַ^m��0b~u�L��~��\r?���O���Azo�׺#��yJ�\õl����f�����=��zk3=C;*ƑXZ-f�Db:��졩��+�@�:>�b���|�QՒ�������.y�Zr��f[ZZ��EmK;��+S]�XJH�zɕ�Ik�~4�x�������s4c=-G��N��@�x��@��2B�T��!�������q�)����[���w��]O���	;z3*���Ze�pq�VE$1�Dc}c����J���I�۱��[�-{�/�`ꗅ�m�V��k�����#�g�/FPX[��H2�D^�6-ml����úTo��~%���P6�V���y���
c��S���ޮ�(D���rԧv���� ,�"�Y�L�t!�MM�u�����\Xk]�'�z�&���=��\���ր�e�=7A0�1�a,��r�EEE]w��MI��+A�^�?b�_�ڬ9��=?�%�����9eewz*�|���H��b��^���6m�nY��������q_ڻͬqD5,ؾ����y�Ԙm�����7�U۟�����B=�Ly�ol��vEo�W����O�O/ع�@wX��a$�`�R� b�_�v�$a4�	wW�
�A��g��ʈ/�c��h���)�~��.-;����Ϋ,T��V�W��\j�f8�5!�������.�7������Wa�n���+�+,cY�x^|��c&���ag��s�dJck�|NO_�Gf��3QQ��LE(�{�3�9ޕ���j���/�
��2��a��ͷ�_e�r1c�����(��U�������P�:_�7I�s�o�#��B��^$xM���"/��| ��,�\~�%�2��0~ͮ�;8��S��M��d�S���%>`U�H�
�FIg��~��3�4��-�eϋ ��آ!�ω"�׸�d��m"��&��`x��%�����S )��,��vD_�1"�q�Y���(��K�YS�h�l���2�e�H�D�ɔE���r�Zƻ�3i*6���'�g�LƻdT6i����D�w(]�w	gl_Gr�>�#^������~�fT$�݃��[o���	�L�����D�n�9��)?�v9�ܐ��098�}�W-j&G@O�ܖV2ϡ礂G(�i5}{��j��B�
[mM�EM��~�����]k�����ѐ���D,�'ǆR䊖�w@���n�D��X�G��J��|.s/]���!2OG�(%l��ݻ�?�N�;�:����:��hg d�Q���8nF�>\��gt�w��
�MN�v-%K�7�����k�I$�Mx��,��̰ᯥB�<З�|�
(J`�<��}X^禦�]�-�_��-L�e�X?�H���*�Jj47��U�8�|d�G\�\���}T�pz�XG�X�J-��ύ��Y�L>��{X�e�-���<g�C����N��ĭ��-�7�*w:�N����W��ZLF�H��U�"<�J���l�ڣ�B�8����hy2%���)��I���*_Uh���&�7`�
/�Uw*]/z�Mp��&�z����pG��ؑ9�")�
:������r F`�X���E��uܑ$�ӂ�|��d�;�D*_����M�V׉#%3�VeM�����ђ�C�R�A�y;/��N:�J�t��_�̚�!'d#*3s$��;��QTV֫�,�]������r�`S9_��w�ؔ�� �@�+BC��r�w�r�&n"��ib,m��ᗮE5��?e��H~�8Dt	}���Ő�7�7hv?gr@y�~����cF��@���&����q�jnK�"�N�!srV�,�h������߿��a9bDjג!��k4��N�k���g�����H���E�Fg�����3��_R�q�H�:-_�?J���AٲJ�XT�u#Yuu�����3)��P�ۡ8���t����KK���D�N�-���!H�r���lz/ŀ�@�}甬���1�B6�~!u���U����UK�m�HW� ���Z|�;�Z���Y�2�����& ��5�����~5=���q?�N�=��ܬZ�)�A���6������,ӆ��i�~��rn�y�Գ�CK�b'<�zl��֋c�;C'�KZ��l����gf�2)�P�?��l+K��'���7LE�쁀^�>���,��B^C��C� �������z!�V���7J�ve�]��]wI#:���#
 �x���XirW��c�;}|�i��ʨ	C��98<|���:~�	jQ����!�dT��?�D�0�+F��J�]��n�|���o��\�L�܏��$v0�����Я���`	����Ya�IbJ��`�)<�g+XA�L��3���Xd`�#k=�%�š��6Y��U��xm�i�Sw�����~�����S��=�d�>ͭȧ��Y`m\#K��ڋ��	ǅ�꛰�f���xhoZ|��7�0��zF�ʷ��s���P�ϯB�j8N���f	O��ln�#��T|>S��|��"''�U�2xP�O��[}٧���m^]�o.��_�s�P�����@ǘ�� �����R��s�\�W?�{����+55"�bOϾ���@$,f=��`q�(�'9�!��L1��+�|�=���0��h���[g�_��_�^fE�J*����؅~Td�188��%�.��^mBf�u�{/ �hg<P�-�\�lv�"�ѣ��^B8���9umh�,ks�(���4y=����:�߅�D�lԬڊM�Ӿ�F,�P����`d˦GQ/�3D��?}ÃKV�P�ؔ�Ɇ����A7���H9ӈ��9��*4����95���d&���������~n��+	s�gw-O���p4�&�Q / ���Ʒ�}Z�vE��OȮ5��n�7�G���z���E�g�S�
\��دݜ�:~��y�o?S��7���i�{�$��������
F�9�P�B���8����3qIIl������!��^%ëOGd�{��{TU���7Wq'�(�w�>��8���HK����T���G�eBzz����ccc2kp���_��Q��O��ܝJ*�h��c���n�U��`����$�[O�)J2^�����햯�5�f5��59�t�^(!�e2@���
(�����Y�=��x�0F�/-�8?�SJ��Q0��������2��f?��)��?=6O��1�����b�_6�(�}#��b�z�N��K	�4w����254�X�pd���/�cӃ���2�PuUW�nD�������:`t��FO���(yy	�#v^�>�{�-�_�5��/~)�8e�3�&�����������c��"_�y����ֽ$�131uO�#\��A�GC�����FeM�,t�r?���䧧G�������w��y��37p3@=ޭ��a&B&_x����J�GJ&���^CJ��Mͬ���l����c�(#������p���=���}2T+����r��rs�i0��Ew��"�i��I���pwu��m�%x������|�hZ�H՘`>l�,r�t-�(i�2��tx�FT $j��Jh	�� |��u���'%m�KH�/���O�|���ֵi���[[�W��c�9[t�  If\􋘷���?�"w�3�|)��OH�����cV�c��c��*%a��%��%�Q��FW�G��}�,c�����;�z��Խ��n��Wk��JԿ���P���_ϊ���h�Z���f��8~�<��*�וBLө�Q?�U����k��]��`G悠���Hˋ�{W�Z���vؔ�jj���?λ��W@����d<(9cc(����u&hM6h��O�_�Ǔ�9�?��j;��>?Y��\�)��~888Ț=��k6�E.5hN ��)�W:���
fA��_p|˭��bgo���
�4����Ʌ��b�H���1n_�O+�Gn0�V�[�01UUTT;��zG����MO/d����i�j�|��P	P%�sZ�͂��EN[%o{���P�v�^�<�ba�m��{��F��������#�0:�����d��KX]`���:^��?�*R�����.��Γ����Pq,L̬HL$�`LqD��)���n��噱�P�x�^�2��wN�y���GG��E��m��"��Pv��k�G�H@��;�G�$������:�dabB���=��|�@0�WGZp(T�C��Z4 ��Ș��$��п��͹����'����˸R�NGP�����L�Of�	d��v89�lT^���X��;98@g�������t-.w���k�����u/.�ᑣ������ڄĬ�	'�gn�a��o���!�S@3��Wc`g72����~,ɿ�Z������{{�j{P���3QQo�So��\���o����fV.n3#%��j���r��i�������GA���d�R�F����o���,�QQNW��3,X����"���)��S�I�z��.��P���X��T��7,��e��h�H��ڷqZ�w�!t�L��:������DTU��JIIٛ���g'�vL%���n7�m[m������nI�մ��Oj4�]���t�y�������Tf���nW ��P�k�^�6��p��6�ϟ���9�8��zwocEbGAf]_!x��|���@�?���m���f�	�?,(��}�4��Q~��l�Q�27�8`/l`�D�D�|��ۯ���i;���������3T��]�_���s1i���n��gr�2u]�h*ȴ�Zy[Ft��M�DM�n����z��>���
RR��!oeS�;�]�ë�E*���!��bMzVVmj��!0�����u��z�5Q��y��g��>?\��KR膊��M��^*�����hK�(�����YYYэ؍j�Z�9TD'͡���	��&V���yyy���[����~K�wI��,,�<2UN�}���j�K�I��?~�k,�궠���{v���{��2u~����s�ٹn��n�p�@'m�G����8��+^mh�#p�����ׄ��?���\A�����ҀyS����X��R��8�����\���t�Y�B"�$ČT
yc���Յ\�mU��ˏN.M	)����O�D�~ǿ���|��������\U�...�`N���LQ�R�K'[�aN��!�w�3!�߅622��e/�Q���A5Q����.]�L"��<��*9l�I��N�.�zl��>2��Z��Y�V�4Ҿ��\����I��k�~����^�d6}�rv�.!%��p��~i���5�����i��esڐLJjې�0l��85,".��ώW�JJ&��ҧ��>�\�Y��Ȝ�˔�h ��dx��[y,T��8Z�� ��8u����|Y��$���TG��ߏ��<#%��k�֥�����@��桥��	l�lL��e���H.ں��A�/FO����0ùG�.{'e�>�2�X�)�">�O��[+�E�K���e�v87?O�Ɔ��P}������A��f�����,��5�:�6K}&�'<$��bz��;����o݂�Fv��]ۛ���6� G��/$ ��WVN��Z.�t�N���N�v�2��J�#�Xxx���7��3H^�G<�"�1 /i7�.��'&�J��{^l����k�V��Z�J���ъ���i)**��)͙��4���Zm�EUKE%p�#��Pú��b�d��;�����AH�v#Q·�]c�yC��ǨS���yN��Rttt�z��:������e���#/��T�Yj�hgk3�[`�lʛ)��L'�����&}MuL�ǣ	���cBtCچhE'����Й����JK{��s?�K����lo�<|�i@��a�������v�]�⹯//+]��x��I?o�ܳ���nD�3G�P���� ���~R&�}��Gp7?���u��u���X8��h^��۷o��iJD��_�.���LM9W��^��3��Cu�~��WP@5N��q�=Y����ـ��Z���	�Y:aQ���G�H'�{�]8>wX�����5kEڣ���H�>��/�g�*����[j����W@�79��*}Xit�����E�����%�}��ihh��,�⨯��� � �]Ū6����f�3��*�[�W�>l9NIk�{��S��Z��M����|V�/Խkln��,����ADB���vD�dd6�+˭]y��O�P�����*���/Pl:x0�`��K��oWϮ����H��^JwWY�Hu�8��R"�����C��100Ш���g�]PQ]�O՟�%)�x�D�3�666RPRBU��IK#�rX!���=��/�S�:'��KJ�\R��9\��bȄ�V����<O��uG�MC����&�sKn��fĚ=w�Q{%Ӻ���q�������k�KH/x��� �B��� ���V/n�2ݼ/��(_B��K�x� U�I�������^k;�D���!���Q�%�y�qqR2!o%G�t�J��$▬���4��ճ��yib��E�e�~a!����{֯�V%kR�4Atss�҇^�������������z��EKk�@�T����'9/�򊾛�� C>��ւ�xf��#.V}���Sذ+7�����{��s��ȣ�_��˳-@fU]�R9�;8�WQ��yn�/]0Qs���魥-Z�X VP-�#�ԝ�.�^���
I�ѩ���̌q?^�``�dݺ�v~<K�5`���=88�<��Ϭ+�a4߉TYє��\i�����afi��W�ͮ�TӪݎ{��g EI\V�%mTTT����Y���"cSS=ǋ��m���w>>>g���reݻ�l3�|�gB�$oQ�KiZ[�_և� ��_��ZX6T���i33+�G��a�tv]H*ԫ�θ����z�4��JA��H�_�TX�iM��p.�)&:��#d7�-�QUU�[n�ed�렴\%���-[��Pq��s����n������bw�<G=ɠjae䂘��+TBU����-n�7��i1��.Z�&//?��H��	���¯QH4)`Tд�S8P����׮�'��,M���-�����4w���Sy?7g�޶fff^�Ue�Z��'P7}&����K��߅m�E�������|5M����!댼Sv J�E1Qe]��z:�
�����@����P��"��˓�a#�	�-E�Z@9?����;һZ�_��J��%���I�ӻ����� �Y1�29΄��т�ݏ1����`���j�Fb3[�I-�?]��"��h>m3�ί��Lp�~�����g鈴�I�l8cb��FƟ4��Z���u�	��)�ggc<c������}	hSn�S�����bg��˺7����"�E34WVۤJ��~���Ȇےt4o�*�(8p�?�/+���9�������А�q-`J@��m�F����7����6�f��`���~���x��[o?�=|޷>�� vXퟨ��}�hl�0c+��þ�~jj*�� ���8":Z:��@�G�ߖ�wt�0Ȅrs�J�f�-7P��� ΰ�@�iwDuu��C�{+<k��_�-��:����ˆ�OZd���d��L}Dlv�CE�~�֭��ֵ�!��j���
��W@T���)�-/0�-���ܘ�j��v8j�юNp����  ��739�fzIa�;!�ɟ���r����j�Q��Pf�n��@�]�I�	���xqơ0O�I�Ƀ�]��v�țټ�GDA�^���6R��֞����o����߈`}�33��q4	?��W ���xXZMG�����`�T���VB�?������zvYI�����P]��g�G�Q��W�skN��� �\vG���]l �N�I�ƪ��Xc�D�!V�j���Z�����r}8+�{iY�g����8Т_,���|��a�P �!����%�PS�������OH@�v9!-?�}�E�%�h�DE���M��*v(6B����Dd<+8�DM�ZVw�p}X��ɜ�<���o!$�FE_#����ݚ͆���ܦgl���ے�QS>�Dhk�v�?��7��Z	�ș�,�:^$Ǎ�$li5 �t��>ط����<2�1�/)(QG�f�X~<�k}� I�?�����3�Zh�.R򲹱1�-����ǀMKlJQ�Xw,+	}�\c-<;<��οw�~� v[���o8���?�qB�����������;Q*/!�7o�e8�Sw��x�p%_�i�iA� p\���`6N��:6��i����(���|�P�Y��fu�4M�v�t���6�|Dȱ����KJ�Q���a�{<m/)[lST���N��&�c^����?�B?4�ࣧ��P��◛Sz�UTx�W�>��w�j�75��""�N�����!�샢�[-�Pߏc�6����jic��`dDf֭�2ݮB/	�����T��C�h�3P��l�p� m1�������255�)$:D�����$�~����D+#�8-oECK��
#�.�`Ƚ��L~����6��������[m-��k-7���:
��**��`�n��O"J��2_�����r�D��O������%Ry�~���8$��L�l�����Z'LRR�����l�v��?��N�IϷ����>A�B!G�1� ������T�a�W�ˎO��E���RQRTd��QB^~RGOoRR[o򣑲�hO���ơ�\�Os��0�����xg�����N�W$��Z���/^�oז���*���Y�i@s���這�orEZn��Xv��֩�T_ׂ�ϯ%�]pH:^ ۾2)�'���4�������V��׿-����jQ$�؝�����##� bh�$j�'q�ȖN���ɰ��ߢ���������`����|�P�w��r���� M�/v7��tբ�A� 6� ���+(�CEE�O�9/p]32I5x����fw��q���$"�D�B^h���	�;t�g5�̕�����cR�������Đ�.���e�"��U���M����r��)*�U���/G��<�HÃf��bW�Q���G+v緢���}��k�}����=dU�hM�@O��ՕKHX�s�L��(0��}Q�j�?�oM��G����3~7Q�V �?d���&O��Mb�4KGU����R���*D񿺗�upS�������f����bE[�]�)ƅf��:�a�W}��'�0h���ţ� Rq�F������@EA!���ݻ��u�>N��%'������	P&B�/��:xԏ�֌'��t`�n6�;z '��q;�&h����p�օ���l_hJHH *����!�X����������"�}}
:߄t�������J���wzf�x]^��d=�nC}l\c��_Ն K���s��_��+Ĺ����8��̱q��k@Y1Ym]n���,�&�J��p
wPDJ��إ��I�D��힁޶(����(�D(�"�q�p��g��^�_���WRR�-�B T��<�&$�*�o�����w�>������K��t������^��e/�������6G�6�
_P���Y��0�jv�Z��⶙��/�� ��)�Z[��>9��\Ʊ�dD�}�j�8��UL����^�[O����w���qzF�75(�����.,�.�e����9�������`���2��)>A���� CH���
���I^��;�ݸvF���z
������*EO�7��Q�:�Z[��8�pfA	,�LJ��o�;Ƈ3e�4��]]ow�''��V'���6)��t�x�PA~X6��ZZ��&��=�b��YZ^��L*�����`��I� ���5�C�������ڸ�ݮO��Ì��{��=GZZ�NL/������J8��S���0)+�pXDjGGGG0q�O�ӛ�!Vz钄��tw?��2����T�x�$ h�\�����\�񴡱*�T��t���D���@��X�������I|N��h�4]߄��1�xD98��̶���{5-X�80k�H>om�wY�2y1. Rֱ=�h���:�ɤUPQQ�o��a0�ZU���~<�d��p�~rG�������0P��E����>6m\�MUF���#M&9��y�S���v.���^������c �l��NB��Ba~GB�~D�7�������^_ ۼ-�ey�����w�_/�f�|:«vF�a����WK��h�O��D@�\g�����w?���-_���)6:�C낭C �������0�(����u~J�X�R�eQ�zI�8,�8R�fs��X�E�X�Avvvw���'K��Q���! Ʃ��[~����FB 3�wTa��5?�#��]�)BW7�mkrllhe�Q�Yr�і��4P�"q?7ٺҷF���5�-���HRA|t�����r!O��|� Y��%��m��zmm��F*��~����T҉����`3����6+݄n���.+���-�!c�W�p�IHxg��T����֓�Vom`%1�Zj�2P�ӨAms�o��`�aoo���o�wbr�`�}TdPI��l~Mc��M����pT_���8���.�~:�ܽ�e^{��^S��6�!��,
��,1g0rH�����������>7&q�7�*sv%6��[}`�����CѰ��C��9�m��қ@3i��O�5��=�{�ܐʰr�^��"�SP@UUUr�G������K&�Z�G�1&qf B�QW[,��"�Rj�G�L�n��uD��LI�� z����c�Z��dGT�Brrr��o�G��ZZ����}�\�N���=���
0��(&9��B��7����u��rW$o{-�a5��̕��op�L�s&"@� ��Bʇj��4쨝�D��*�v��QB�풎��&I؛�L�ޅX$3FD؀�ړ`��f����놺���_���z�;(��9vף9�'V@�׻ÆZ���.nuu�4A���nVÞ���~%'!>�:K�"P<�^䍚���vNCm	gb�H�����Lm��P,,4��
����bA���t�50����>8��� ����������_���Y+�
�o?��l$e8ڛ��6H�_\D8Qr!��T[ϖh��{�jii9ǐ����mvm�Ɖ����������-�W,��|��'##k�v���` �[Ǿ��t�,�U2_I~B�����b��_KHA�|�F��4�v��.��btp9,p�A�G�F�_ºr�14�&@���֊,�������V3���Y-�;�����cv�.��R��8""�7SSi=��X
��z���2���9/}�𐊏���?��?�Ft��&NY�������|�]W���+)R��uc�GI����t9��������Ț��@�ZB�K��O$��@M��/$?ѯ�����M�qM�Ғ>22r�$�Z>�%$3��ĝ��4!�O%*��?[ESµ�nOQ���#h-;b^�H��:���	�I��'&��ka�ID|M�"U3�hmDlYyy��r��zF)� ���+���O�Y�*�$&���y�����H(�J_RBiݡ �҇W!P�2��E�G5AM��E�o�'��u��~�xkw�ƺ 77���LW��F�>5s�|N��*��6$�y����G�|�eϠ��u��������������?����kGG�KU��/\��ӳ����k���z~�PV��m���<?�f��y�,���aVSS�3!J��	L���21I��C��h"���ML ��'!a�Xϗ'�r��h�X�*�EՊ���c��Қ@�n�LO/Si?����%�������\Wtૠ��!����*o���e�0�����2��Oq�c��a�����::�==�B�.`���$)
�[D����&9���|��ؘ��-.��l(ؗ@0!##��a�;��������7~2a/j�"@i_���?03��g����
�<=�y��;^�7�Ԃ�x)`Ɗ�$B�B�Q]]ݳ��n�Z��	�rZ�Hzz��)��;[Z��v�qj���lp�E4�EĲ~��>61�����g�8{��52��{ǁ{ #�j[�h��}�ݍ١*kD���̏�xN��35���ѼsU^EET�b�QE����=��H�n�#��!m��VV?޾3��r��eY8���Y�l?�4b�/��&���.ܗ�g\VV֣�z壹�tAv��M�޽3�[�a��5�I�d�X�R]]=��f��k�h�%;BA�WoO��������j�Z!�M��Wp@+����p����a!!�@�3� `A���m��{��v������\�Ӧ��ݹr��9��|ѡ����) *L���~���`�TLʿ,�UU���a���Q�}����;��bkK�����k�Q�Q=��(^�wɃCC��c�/Up����**��L\�ޛ*R��6���<�|�|k���������@��|Eb\||F�ݑt�8�:T`U8��OOo�����J�"!%��� �����)� ݠt�HJHwwH��twHw׳���~~s]��gv�u�׽�>g�����Y��atFۯ%E%�_��R�#u�Y�|vv��n�s0�Z}F���˸�����T��%��ZSX8�	,��x樗1cP�D��'&jZ7��1zL��4�p5/=�x��YO�Z�����Ye'f`�S�|xdd�+��@P����G�L��9���^���<���?�&v\�x��P�g[#V�U���ɲ-k�����_�[Gmi���Z�~d򹁺<��|���~��fɢ��z�K3\L~0vPJ^���lL
���K��{��c��&���g��jH��8n���%SF6
Ap��Of�sĤ�pi����?�}N'� ��`����@�:J���!�F�օ���h�O��X�s5���J@4�1-X�<���N�ѩ�'�F���!����l��V����*EF7�t?�t�_�RKE�?K̚�t�u�j	�h�<�%{�߽��6���.���r����y�f��M��߸==\��pTv9Rd�l�䆭/����~�u�{�� {�U���Uwy�>S+  �5�N$/m;�����)���C���d��H�!�Jl��p���9��D�c�ޫ�=��^�r��3��>���>�X���g0j�~��?2:�������SR���ݮ���?��1 ~ԁx5�O�;�pK%�ioo��w�d��b\���uc��P�㮑�Y_����:��J�Ub����ˋ�K|RRƂ��́<mj��m����P���6r����Ůhy:}���?F^mt09�0�^�Ȅ�����#??{���������[��[n��4�y�>O�v�l���x�)��EFG�T;���"D�yw���nM�{n�Ԝ87�[�-���N��Qcn��~�%LCԠ5��S���{U�c<&����`�����ÍH����R��M<�8�2^M����/�`U�GO!����`�,�W�,&\�1��WM��
Mp;�e3�:?�upp�t���x�d��\�VAA��RB�\Ol�o�{̥䕗ǖ�Q�q����3�ݎ���1�|}�?0J2lL�|�@툎�nko �cnL�PM���]ō1�w�u��hxyUy������=���
�k��B[�����{�M��m�3�JD�ώ2�:�ڐ%0d%��Z ��++]]������� ��Go�~��Bٸ5�^8��*���(wyU���f@����eo�ܿ�eף�&"dM~a�yW%�!W��[i1��� �Ӄ���xb-r_���>:��H&����R=�%���yw�Oj��xeI�������.��?�'d�E3 ��c�TW<Q0�����)���z(��[[J�q���(;Ԣ�-/�<���a��j��N�� APS0�YnE��`�IƷ;��1Ɵff��m�)t�[����
e��|w���eJl��x��
 Y�]GGO|���c��I�/��3�5�HV�?Վ���"�s �bk�)))zbJ����%fd/�o�r`ݽ�����5<�2���������z��"ǲ�r������DO��_$=��L�0�z����|9gj�f���M��������������a��>��x�	J�L�P����Wݍ�*_j�#40?�Nb���>�����?~��>~��f���$������۽�=�������� )�l������_������:�V@������N8U����i"T����|�NҔ �ɂ��VP�L�I汱��3��������ɻ3������+���L
���WH �]O�2�����Q `^��J�*��-]0	�i�������2��ˌ#*�Yh&���e{��e����!5�ӷ�S5@	wd;g�rP��b�w��Vr������� -v�W�[�_4�[-t� �- ����yc4LLP"�����W��s�|��[I��<kYG�K}͜�y��i,�m�9�9l���S7���&��g;Zb����3jYYYӢ���ځ����N'[s�l�#, ��J�0���6m�+J\���@�JZ_�4<D�m�R��Ll:�H�����^�l[wwDF^@ v��3)�}#��|�!ւ���|�C����b�^�&\"���N�,,8����c�ff��٪Gs���F�7oq^�ƴ�
���fǚ�<��|uf���d��{@�N[M-���qv�d�E�\�..�d����<]<�:���\p���QA��<�౫��a�;�):�=��;Y^�o�vv����1JEm���Y�ۮ*yO���C����G�a�_+/���K3�����)=�I�[�ڳ�>a@N%��`��-�+��V3�ζ�>$ໄ}�����Į���8x�G����+��Sd;����3�^uQa�֜�&����	7�)�Cʈ�IņY5�=���e���>���Z����]�>vKz���ǘ�rV��B�3����۷����g8d�
&��_9��w��o�:�L��
>�r+h��D���z�WO=�:��l5ߤ�t�9��&����P���1ja� V��ׅ�������O�oZ�������i��f�R0�X���+��.����H��k��2�X�Ap/�VJ�RnVV��J�GJ�gg�\���߮	f���`��|,�S�Z����ŵa�Z�2���୐E�ϟi�ƛ��jiia�v�@(�-{�}tr"q�c5עRe�Ӡt�{e�t���K/����J��;��N�=����+��ђj�c�����S�e�^�|�'�,Î����>+��KBE��`��7������Y7S\�f(w�GZu�{���� H�J�i���ď�E������l'P��zxx�J��u<�l�����84%��,,�����!�Pj`�$>�>XWO�CN�C1�ce�	��И2;ˉ�ʯ���w�(7uwb�_ʈ_+�Cc#VB0Ƙm����ak}�n���ׅ5 q���}q/ood��KY��Q�8�"0�?�	�fR<��^�K�k�CII�Շ����p d{ze ��a`(�R^j]�$Z�Pq��Q|X�r�b��c���J�@�����X`���w*�����AEx��鑴����b��t�7�������O��ƦXXY[zS$BB)��^�%��x?)pG����{.���Uv��+�s�HM���=J,W9+�X)"�X��}(��ϟ��3�d�5`2�Ky��oT/B���n����lig�T��_��k=Cu�'��,|���n9��^-%�Ǎu[M;����J[�ZW0�&��cuS�O�׮r�o�ex)%մYw�jG�H��]+���};�l���1�S�8L�B%4>�ʿ�)w>�Ů[Ŧ}��d���JKK����>|�D/����}j@>=�]J��"Kg��h{�|Kؒ
��0�<ބk�Z���Y�U����O�T��V]B�2����9=g�~�:�A@'&&�����ܤ���7�����G@��~�2J,���`����נ�/t��,�mn�v~Q�V��1e��jV4<H�m��w7�r'x`�����P�#���|�/�����Y���%g&����AW�~�V���PN��|Tavb�x���#�sSeee33��<P	^����b{�Xl��!�	�4eby�PL��"���S-A��+c3�
�`��� �^��-2y��	Y��C/��س�� u��FB���+�!#���ab/���|+3��"�s-�K���=�w���9d�"7^��>��\`9�;��.��'��b^*-.n�T����:�NRb�����ip��Cy,9�ך��1=추8�5�	Q{��:�x/ã���$��=Xu27k�h��%�h��G��RSS��U�u�>xQ�������_I�]��u��`�.����x$ֲ�ް]��A���ZA��c��<)-KJ��Z[�}�FB�E;f�ne�������ߞm��Z�y�f�x���'����1_�e�w�?������?��D��#�����w7������UW�(�V���b}̻_544�Tٿ/Ї	W)6�"'le�r�B	�ړ�]fA�"�*���h���P��xS�蠍���k�e��h.����;bb~l۫�6�D�!zH��&'K�ǧ�X��FC#H,�t�A��P�i[��n��� �)��㦟t�����Hm7Յp1Q;`d"B��ܶ�p���ظ�/���q�C �������ο"����������Z�G�B�?7����,���^�<ad�3��ٵO�ϸ�����x0��_������խ�����B�/���kW~�,�(V�+[��&���upr
8�Q���~�@%�G����	]��(��h�蕶������G`Z��������u:8;s����N�@w�l���V`f�>�]h�7��P�!�]��yNb0��[�z0ꖤ�*Gs�����މ����E3V��u�
7�A~�iQa�33s�	��Y��9'g�(		���BG8�v�i�;��9Å���+���_��%�g|�(���kƋ0/�x�
O�k&N.�h:�v0���ДH��D��c``�E�ڮJ��F��A��I����N����y�/��E���_w[�K�\^^�n?������2��&k��&�C@Bm���o�����=���R�\�4dZ��qX�8?%�oۥ��Y���;p�{���`ìt����"�|Q�C��%�...�Ty`�9��u�1\,.-�2�B�H�m�N�,DDD�C�ջ�љ3RQQq�
޻�;�lW��z_o���4.�:�uK���a9ڴ���_���)�X�y��=1����A���/����pqV��z��7��ެ��rI�D1��D8��>�y1�G�[XT����tV�����G��|�n����O����'���{��`��f����O�l���/��Y�fnV�����
J����4#����:�q��}�TH⤖��\j����-1��%,���Q+�Z�n+U���V#�X >��׉I/3V����[`2R��m(QE w��c*j]O%����B�C�r��-�����a����(��4'%50<��z���)�:���z���]��bY��vXUN~����]�5+��.�-����IȞ:��D����?^G�}���&����D��]�dlQSn��}\�+���Fq���H9::O.qpp}�N�TV�K,��C�^�D���XV���&��}`�hc���37=F
�}�� ����̢����I�#�d%��		yCW���4��:6�qs�hSm���� e�h;�{�@��߯@��Ǝk}~b�긻���˞��̟C�֥�2
`�>P�-


���n�9o�Q�o���D]�~]��B$�_��MC\@fG�ncTy9���w����_�~u5�-\�PS� ��M�LH���i}�z��½t�#(�g���S?lrz�:&�������2����i�ܛr�"r��.ѧ4�=��wq�:Y6��h��ڋ�X!��ȹ�OQ>������j��s����j��F�@��H���^���N�paez]�qq��^m�NHOO�G����oB�8��=��䬊�=Ɨ6q&b=�|̫z��vk~)����?���Β��J����X���u(����[������؈nddtG4MC6^���0���s����Ǥp�����0�"/ЇP��m����9 R�V�S���[����5��dc��d����ˁ���鵵 �Έ�?~�h�30М�&��hK�gZ������JV����:�\���&r6�;��������`Ɉ@E�<F&&LPIJ.//oi�"�dr�,���m/�����J��@N����3~��೚���BK{���X^���^.�o#Վ\�g����Pл7��~��j��K^U��]���oц1���������gY��������,5������S��b�b|�+��Q㒵ר���3�-�����Pju0'k][Ӹ����^��nj<f�/^�pc#����v;�^����UnƵGu͵�2�X�چW��0��F�τ��/R���]^�/�VdJJwYbdj����|1*��IRQU娲ߌ8�P	��FA��@����[�G��E(�t�����A�YY�F\��ۉ���=c�0�$8=i�ڱ6�O����>Tk���Z�^�	
�e���R-4��+1S�y���� ���g4�!���jgSSS�ާp�I�Pмb��wO笙�X5�.Y��ɑ;��@'$�zb��}b$��u\\]V%Ύ��_7�a��H�lZMq���m�ߤ�D$��v5�ɼĬD�3ݬa����^PS��C�����Z�8ӹ<hb��?����HA����g1�@�b�� 4�p_�,(����ݸ�:�ǵ\\�腺���V��T�TT�x�D��WvI�����Z�||$0�b��'%'G?T/e'b���.��30h*���`Q�֑I�=??�~�漿B2���pw��N�(J���zI�ˏ�fD�iwg���L|�������ٳ.���� *�����md���	� F���յ[m�v�Z��c�/~X7o^�5+�F?2�ڤ_���J�X(��Z�y�՜J��0,{t�O��A�eT��;�����(��75�Q$VEz�L��g�%���c��A_�Û���B(%��풪��7)��~$al�*� �8K��R�Eǀ�ڸS�U�m�&>:��j��g�˃&?�ƪY�r���)ga�j��Abh��6�9`?nh����.2����0}] 2 \\XXX�Z�9�]gǻ�())�X���n{�SJ���l��'��(/'7����c�h���!�t1�q�r#�V��d���O�j�cB� 䌯�iaa�縸�����%t����`������-�ꪵ�u�����ߏL{�S<�w����癃�R���?�BɁ��>}	�+%MOK�W�n�V�Դ/��\jU��7���Q�f��Z՘T��3G[3��+
wx-=�afP �! ��P$Sm��@�B�K9�e�������]0'|y�%��[<��~]��>��Uk|���t��A�ևP��C|�WU=��/M`dd�p�d���@:���	�!�;�6o.��XY��.Y?ؘ����+з^���7Y��v�K����t(�v��euvd���kM|��@��.���w�{���jn�8*9⦦��)��,R�i�໴e d��ѡ�������q8��a�\^Y���l$oiia����}���:7��Ցa?88���=b�+���d0OO[[�[D�J�$T���Ͷ4^���Q2��E�����-cc�)�_�.	0�v*�266�N�Ip���j����*�����߬���ipnh���p�Ԝpwg�\]}�y�מY��0�0/9��aX0�j�a�Ur���"���)�vX�B�*�=�?6��('�����.0���?�7�
_���"�ۧ�3�6]�V1�R\R�0�� ���#%!����eS񻑯��*�)��Py�TE����ފ�����\�����!쑕۝������trr�&3x���y�O���j�G�N~C�b�S!R����d �����Δ���11���ii�,9P	�uپL���8����*,�|iy��U��ӧ��r��u�T���z�RRR���!��?7�͊�A���a�y����R��'��=-���kk>?/������'����f����M~�`��\��%%%���s�;k��I��G`��E���\�C�c{�:l��
��H��o3��vt �� T�o��Swf{kgG<y�ݺZI�Dzn�����Pj�{���������_Eh~�xK�0>���q���F3��
@�����b�9��Cnc�uRRr6��˚��/���,%���%�{���d���܂A�V�.��"�������%��c�A�#5k�/2|���3����t���f�~��˳�����P�f�[#e��af�>zD��k�zc1���iמ��H _4vvJz�u���:����6(�69Y��"��'G)��c�9���(!�'���D��������D�*R�
��p�-�h�y �3fxx��/�]>���������0�YP����[�>āj���x9�X]S���F�dgg��2U����1��?�������?����w�����,*]�R��Adl��7W;�6�����^�Ӯ[d�y[���?�M_������Z9�o�]Q�zS:}�GGG�G|<��
���&��<�k�ٲ�ѡ�����2+�q^��y����	����sLL�����'�%%�h�M!��:g��-�LL۾��cb�z�z{���g�B|�Z聕m��mI���	��B�"�1�ֆ=s��W�3��ŤN�>g���7���a�Q��z�54��m_4JW~��se:����[S�D�RN�@�2WO����c�Z"�6���=���s�_�������Wڮ�[��ʶ�ҢJ��g�4���21��緗y��ֈ�Vg�&n#{�r��D(�Ϲ�fy�7���U��/�x��^e�u���v����q����W�\�����4C�)1�l2��%7��Hx��=���Q�ׯ����yZ��N�o"��Z^De$���8<l�}%)fR�~J���؇?|Tmo?z{�� .�A�N�yk�H���VYO��T^�o����<������G�&cӲ<��R
@�S�5$G�����t����/^\ONIax#@�JZ�$kuu��<S
@��~��_�8A�����7�4�N���C���f6](3Z� ��M*W<=L�J�}���XF�#�@����ߴZL<��TS��:v'S����chq؞����
��4I��vپ��,M��8�ƾ���89��z�K���"��ɩ�({qy�!����|�H}'���~?��tg{vv��ӷ1�-o3MQi�?�V5m~���*�P�o�k��8�ݏ{D�x�KE��^#�s�8�
��D�n��Q��	�<g����qA�ͥ���f2���Ļ�RR�&�Vs�������(~*�T��q��Kו��a^�B���<��?}��rx۠�0�,�[�Q�&S���'}	��zڃ���Ζ�����yޑ2� Lg+Ys�MX�Գn_�!��"I��I��lm=;n���Ώ����0�ƛ�52���MIٙ�ũm�]O��Hh嬃os����L`�����{�`��.(�ww�����Aq�^�e��������t���S�$��5pL��X�"��+�d��p���\�N�e��}oB�w�7z#2!A$�-�G��)!����l�� |�+?f?c����L�[��t�bS}�h;�wm	��Z�ɳׯ�?a�!�los*��w�j\R����_`�����-*�|�-+ߚ���g��������/���3I[��2�Hʲ�0˫i��X/�Я���V)������Fw����FU��`��<�Ll[�X����;)))R1���1n�Ij~O�2�z8�ܼ�~6G=�`��{p�fՓ�¢">��|�[����c��D������Hލ��5̉Ʒܙ%bU���z�����k���;��Y���=٪E;N��%�^�"ϟ# ��P �Zh9#r�Y��r�������'*��خ*��O�	���v���H��Mh������������|�����	���?�TR��{ܟRO?�6��{�T�H	^ F#�C�hy�R��ޠ!�;|���_����(s�Ŕ�꣛24�����4[o�Hf4�"O;�`�tz���94G>UJL���]_��ϑ'������`N��_���3?�ORv���0Ǥˮ���`��4��.��96p��CV����<4�����ř#H�U�jnrd��^��%[ݖ ���~��L�����������ѶL�ޞē�w|Mu5�c�ؾ��BCIF���lB
9���5@�w���g�u��֤���cy�>ݓ�6첚S��Ո�_4�0��/Ҷ��3���|��@�?  ��i�0�(�<�+��L�\ˮ��Ѽm�׾���]����C!A��򳳳�Fꋧ&&L���������;]�����u�e�N���:ȁ��P<OOϮ�@@U�1���[��|�i� @.�B��]��IMFL�o1QI��
��{�9PsP�V��O#-�E�Rcy���^�y�;��s��5��P� n�ޟ2�˓5��~�b�*ʽJZ�a?庴W�*��h�1���<����c��m�	�R�>F7�j�CǓ�4̀7��]��]ζ[Y����M����e�|�ٰ(oP{q;�˸qq�
��0�������a���[�K	aQQ*nVQ$��|�'��`�J��F �R�L���.���=Q{�s%=^����r�u��{�����\@:|�x�a�%�r5�s(���lV����G�CoR>�S��Vfqã��q0E�%Q[{{�ϟ^��z�}}�z��Y���f!���i	`c�/���`}��[���Q0G�ȬT˶���D����!��Vj���s�*�g�%�����
:����	�z������K��4�_�,���d��%t�����m�C�����H<\Qi�_Y�m/�5��q��hǠ��,>�Z�eB�����!3�ó�Pw��ߡ�M�h���-��_��,Ӫ�l������_pp���,�Π_�0�s��A��6k�t�hY>d�㋞�7 빹W=&����)r��L��E�f�]���Ɍ��r+��G�rZ�j��h�������v��̑D[�/2�qR\k~�,u3�O����4�`^��|���.�Z�;SG���fA��MK����%;�.����uJ��	�Y��������]}Yhff�5�r�vHs�I�o#.			fMn7�Z����fG#�#�ⲳ w�R.�'psrrj��U�ob"ָ�v@�B��Fa�(��h{.��ڮy�8�M�vo����6�|�1��7n��>ONM�2��u�8T�������X�ہ�S$	[ǭ{_�v�5sV�v�k����Y��� �\��q��?6K*}�����t��,q�Zn��i�_a���ҽ?��u��+�6�ճ��������d��o�" v�I���
�?m�Z�-DV(K�e�����rx��Aw3ݷ��/_�<ss��x)Xd�Iڝ �}1<6�]����~oI�)�f�U��:�eTL굂B�|;���`L�))_����Vwy�9���n6��#�-]6J�@�����r�z�;�Ůh֩1xdr1����Q��c烵��_2K�����nw�2=2�lQ6�W���Q���r���� �PG��Ҿ��u�W�u�V�'�AA����OHd(�'6,�E��K��|n{���G�D�K��[y�4F�xCͻ�B'k=N��;!����i�z,ʸ �#�Z�������M?<����r\]]���=���a�� +�~�SR��¢�3�n;������E(��LŬ��^� �?�$e�~�6~%�~r$�u�L����vW����7��N��9NՄT���2�*����$�IL�o�	l��w��g�-���<�B��Oq������cށ|BaB���`���g�"�.��ܹ��gߵ��������{R�
E�fK��s*zo��~�d�.������x0 ���l>��ib����5N%��Ѭ��	�a��̆X�.~�~8W�Ӓ$}�����ޘ�*�D����>�[��իX~�H7W�R��,2<�#��>�VU~3�ȗ��H��_j|���t���ؓ�~���tl�a%#-�"j����������os���{�IXn��Z�]]�i�z����Ň+�%fC�&iK-&&,�Z���>��-6m��x�k�l��,a�YJ��G��Q��K�%f��\�~��p��X��HA�����SQm��f�����<;7���[]Z)&&|瓟Ϟvԟ!��}�}��fU##ƾ4ټ}<7QQ����DG�+��M�=�U��$�'?.//�>�ծ�,�S�h<��p�8�v7ڷ�S^ˡׄ9������L�ryy�88�ߺ��j��&��>Xd�E�8��'��V�,jO��I��n�%���K�\702��N5��g�EBFF�����Ě�ʅۈ���qη9V�7�!r��x�ך�-�!K+�.�K\�o��ϋ�!�:W{��i�a����J�n���Tj]��������-C�Q<���I�yܪ�*Lo��<�r5@�L����h&kID���(6����*q!/s�����?75��-
8l�@��&�������R⒳{0HF(T��D;���������E�+���N��I��Z�RK����r�~�;��|1H6ld���S���1:�'U=m1輪9�kE=m��v�i��JNU�i�@:U>Tk���F��fuXll�L�!�_L<�4�2��x�*��W|ng�֋]On � ���I%�O@�fI?��h���`��_��{{{1qpn�g`���HIME"�Tp�ˋs���^X�6}�29�e���?���}�e�[�����J}����H��K��Ɋ�!'��%�~$��53�~�����:?SF����OV���#�=<�"�ӛ��g��� ==�ו���/(�&@�泲��DU�-.#��	{�fd�C~���/�JP��KL��=B���m_�&�z��T����|������_H��T�+���#���O�!��v�waP�)�'��y�wzGHIz2���5&F��~P2c%�U�А20��v�# �7Y\�?�B-$$dq���1�.ŦD��:�}�q�n
���N����/��ڷ��}$�./벸����/���.��:�yM&��ED��U�e���#�H�kp�vcH{�����O��(�t�uF�٫��O�=��{���Y��c����_�롶��w@b��Ο<����[Z���_Z
�����!˖�Ѐ��$c4�K��9���܃��/������u��QsE�͌iV�"4��d�{��{ɉ7��=��Ȉ������~�ry�FF���z��抗�)"�
�l[��h&Z�����[��d�c�5�O�*��SF������˨�
ڃ��걁�$�N���l�C�����5�*Z>��5�~�z�q���
���=�N��[L 
{Cχ�>���Z�ʸ�)��kOx��5�����9:�����+ɖ�Ӿ��9�����O���x�k�	�+�wۦ7�W�Y����]�-p��7�w^��Pf�(XFR�p�c�l�y�����1P�b���3��Y��k�"t?�C"��}EQ(�)r��'�{I.���lV�6��=�G�i�+ׯ�iR�E����#�47�/�PLE�����J�Z�2ӹ���V����}����۟�Z��ׇ*12���7��N��Q�3�B��+9Z������"v,����:*�Z��Y�=�&:��}1�;����,��jR����&+���Q�8՘,[X8���t����y�\#��G�j/�{͇�hƬ���y/s���З�Fx���0�^�Ɉ��|�� PK   ���XP��/�  ǽ  /   images/f42d805d-3c79-4d19-85d7-77e6ec425ca7.png\�T����"  "%�R"��%�]�J7�ҝRҭtww�tI���<��]wݽ�Y.����;o<����U�GA�C���A��Q���u��y���s}X��y�($����������H����,{;)�z0�VP,~gN��,khm�l*S�6f��}D!3ܤ��VR�q{�Y\ÑV�]'A���fӵ4�ϓ��q�K����y���q�=~<I�����ӗ!hG{��%�M?�ă���w-&O���;z+8��Q���f���~O�&��D���?��e�yJ�@�-B�����z%1�����>&]���b��bp��W�	�H(a�o��d��-���Q�+4�R\�xWe���*.4�����oq�`��F8��c�L{p��ڢ��}
sR��z�S�!�����w�
^~&�*]��R�\H��sݐq�g�A�*�{��p���_���tcd�=㬖T[`��e�b�^Y0>Y��҆�R�L���y��up������$:�+􇇇�q2o��h�ۮ|�6 +ݐ����%T��0+�U����"���7��\��A����'��KF�R���������Jy ��a��υ�;�f��J;��	}|��j�b�i�]�|$1�\��s� i��~b�ͤ=,
�Ȁ��I>��[$�m��-"�c�V��g�~���'�����K��k>:,��.�"C����H��3�_$2^.<�U��)�	W����
ٟ?���*ȥI��+̕b����b�
�Tm&��J�](H��7{���w�xc��%"ҽ�Q�Ύ���<���Ͳ��kNtttfף%���qj�ES���.���8��a���A�Oԧ	�XH�?�����K���s� ȸ4w0��.��\�g�?��涉�Ȃ�E�L��/ڿ�q��1�w�0��ßj0�������@*����8�����E{gm�R���AY%ߣ���<,�QO}�o���04��=����_/��W��"BB�N�l��0�\@0~�h�U&H$�=��?�W��� u���YLAL$��Sh�,�٩�ha4b>�<P%oɁ�@����S����ez�R��M�/6��C�i.f�����oӳ�������S�ae*���r�|%�|%�MV��0"u�T����B�l���2w�$����u?I.�ꟆU�nn80�����00x��0�������CnbȚ	3y�6��7P�_,��
D*��{y��?�%���&PRVN�!��d-O��6�_d�����ѫD��,��V��c�݃�k˩�$^����96�
Ll_Q��z���)�����%��'.�7�ٓ����>�$g�_�1vm����
	B�^��z�t	
��;"$��UU����.���f�B�փ.��'�����뙓 �vHOW��3� ��S/
�����?vW7��KF<jF��Z�G��p�����V��GF�;�uu-7K�Ɉ�(!�a]�"���T�OM��<7�DE�待6���V�!�iJ�%9�f��f�����S�?2ޤ��CNS��m��^�?=�b��vjwZe����R>(���/�%�SF�'�g��a��渶�0n�C6�l���_����o���ͽX"%ُ�
����cka��,x�|t�|rE)Q���;��Ի�I��_[���W1Նp���eK�w5���b��k!0TW;O�/:"��M���{c�;�_�|E$��E���+�eE���K�k6��	+7�-��I�t�S
�^�r#^���Hw�k�����!��#�#�k�K%%�<\����D-���M�=	�F�dq�8�455[|�$��42�˖�p���c�٢Q��X^E��\�:��祺���Ĩ�sh��7n���sj���i(2T�E*aY���;�����LoD�Ă��G�����=S'owk���K-x_����>I�����D���Z���Ͽj9��!CO�7���{�K���dvu�o�W��aA�sbaqS)�1K�"�w�Q�ӳ���,}9*�΀���4[(���8��`��}�慀!.�?�XT==��0�*T6Ư�"�ڃΏ[���l%E�R'fH�p���E�� 4a������ײ�|�b1�c����aID��9wf��X��Ku�0���d�0��,^�c?_*��+l"�.�������k���Թ����ܽG
u.6%��M���
br��O$�N�?�?�bi���ܛ�\~�u1t`�0�AS=���~��3��e>z�����������uR�@�h�|Y�+�9�qM47��B���F8��&��O���\�p�}����uJ�y�H�k82z��_��9�"�5��`-��|&r�LS�Q��+%BŠrV,*����#om�.ל� W,�}9�@�p�H�����'����P�6�"z�6���?����aF#3��|8��?N�~{��;6��K���14��p��% ���8[r��N�Ȧ�B/��W)���e��ckm����"6I��ߺhwFDD�WEB��(qM$2)�X��E�/��$j?0T:9�TU��0�||��M��sC����(e����jZxU׷Q�
�}��i����D�۩a�� p��	�SvG�'<��ƾ�ãV����	MM︤е��Xp>��%G���*ӕo�"]�b���Õ�P��el�{Ԙ�� @2}�HI�X֦����ݱ11~7�;w�����YR���q�����&�����hn��,��Fg�؇V�S�^���>��.���4�榤}��������Ot�"+~j����"�%�`����W�
}m�?eT���u͝�_�Z&L�F��CDL�����9A*pkkˏq�pq�⡮���?�xW�I�v�SR�S:���J R�U��0�-�u�T��!c\�W@;Gj�p�Ic�tdd^��6��H?�v���_c����Q�C�� _��\mh�,,ts=��D=�T��_��+���_+��1��"�.5Vѩ�0�9�HW�
������NŰiL]��㝳��ԓ߆T�b-N4�X�!�ѥ�*7 N8h��׹��:���0�OOˤ�_EtَD�b��ţ|b'�
ޞ���QȐc�7�bq�b2_Ǡ1Nhc�1Kp�,�P�Ģ���o���F��� R��r�eU���mWa���Ƨ"�9��+k��uZ$�*6�Ud��Y�̪�a���W��b���K���t�<iק�)Y2�p����Z{[l���;=R�Kţ;|6��x�Â>��&�h��L]Q��ȒQ��W��\�E�����8>�A�����,`�E�� �y��7����YQ,�˧6&~qk/^���m�(�M�X��O������_�.s�E��L�n��PBv�l#����c��J�&�<������,������>ߧY%t���T�>�K������&t9
��چnA;���	����"����?]p+��hm!]��r�?_I@9u��g
G��\#��Z:O��0����5V?_|H��
v�x�&j�\ϥ�W~��s���z�ֻ�!����	Ve[�Su��梦���{����z��l���kr�V���s:����G�M,�<t����ю�a<`%
�g8�/�lG���'���n��.���y�y�0@�Ȇ|A��[���_cbR��"�pj�;�=iD��YN�Uv�����a|?<��1�+���ĥCA-�c�ig������D�DDV1�-���DMArѿ�_�m*���������²1X�M����X�t_����05��0~Ã��<��m�=;�M|�1y���ъ��݇fB���f�R%�Ye��4�i�S#�I�{�y��{���ȗw�#3U��~�#&���ԉ�ls�S�����Jb!v�Ϋڨd�{|��a��b<���0
��o���ajb������n��
K��gr8_f��/<��W|���V��20�"O5�T!6i[m��Yk|�Jhy���H!x�%�A1|*�v�C���h�h|j޿U>��Z���'��[��v+�bnv��@S����Q.J|<Mn�";�o��Y�|�[�o�h&ȩU��Tc�p,p�Z��ҼS9|�B�e�:=S�e�o^|�Or:;;v��I^��K�5^����.�͐�ު`�p����E>�á	E^�a���0~7�A}�e5�����.��\�dHu�3����ol��b����1tl��I��?��ҿc�ś�BQ�1(����"Y(��W�����=�z���7�Y��mN_5{�z�,
&�������9�\��і���-1$�ez�M�o���E��{�֎Kߞ��b��s$�J4�v�?=ɀ�N�:���Ԋh�J����Ս>N)�CJ�FW�%���iq�t�0/Z����0��X_b�ǂ��4����S��J(DG1ĭz��.-��ѧk�qpK(1Q����q�]X	�"�C��vf���*�Dy�`�����ǳ�!�-ň���C�/oq`��Ia��f�K��4�s�:�^7a:"���\�+{g���j�G�3z��A��+?������h��M(C��v��[�NP-&���{�e��O���q�!�9���>��>4�WX	*I7�;��݆���V�5��� H�*N��zB�I��}�Z��*�n�ӣ^fk��22�;�iqf���O�n�%����$B_&��W�������V>���o�Ҡb�W�&Xߙ6+I�RM(w�(A�`'}7���t+�sC;���x�������.S7R����eQ��f�&('�
�� J�&����FM
< ����U,|Θ�JM�_;�p;�;���N_�^T֩K�b�{AU��6�1�.5W|�����|��WX?��՗�|�N��y�lyk�V�����w���H�&��W����VS6C�+_F�}���5�ɪ>m'�Uźi��9X:(rJ)�����w?��Qu��!>T6�.�DsTr.jvt�|���k�C����\���r��~v����.�B�� �G�i�xJG��˗<3�vv�F�A�B賜a"Ga�_��ε4c��ɽ�:6�W�M�˵��B9�q������~=M�n��8�a���������[�P��
���uh�����A���g��vF��zk�/[��aM�������L�sR�ӏ�Rԯf�T0wE�3�Ԣ'�jl�;�0ˊ�=�6�3AuH��������0�7��F���XKX|E9#).'��FK��
װ}S���nǂ��,��jo`�Q��l+*�f�N��ox��x<U�����Y'��2�P��sɄ*��]SַHf�t_�!ى"B+ђ� t*� ����W������7p�_K�UU��Ⱦ;
�<MWZ�1�r�'���$��R�E����1D�C=�Yi1����U���_nC���	�d޲��?�h���:6�QJ8�vB`Y�CjP'8�̋���%�D<��2	������:V�`��<�#�<��P<uK!�$�Ԍ-��ѫ��@>@�v:��Z��n���a�̆ONl�_|��Ϭe�2��BX2Spn	z8H�P:��r��N@C/V;�R��9-S���|�W����*	�m���
��9���!�^<E��#9�%�!�qn�Ÿ6&�4zU]7K�yQ0��ͱ��?n}^�WW3O,�K���7&"�S�#�>�«���p6�LN���/�2Ďywtq���$x���S�������zh���@�ʾ��Ef�S�Wt��z�e�A䳴h��F��*���a�)(��
�
�mT&��M�o왧8������n�Aɍ8{M�6�Y[�u�Oq�ᵃ�A�׌�ڴ��RMK�-I��m���ϘõdT[��SW����t���*N�-�ҋϲ;��%	ג741[�y��h�"N�,�_P󣄗�V`:��hS�xQ����j�k9��3bCHԓ�{Oi��#{��dm�O��	N�<�m59զb��#"����ܵ�q�[g�x>�M66��ZC�h6��?]�K�X��c��ta�p4{Le1e�i3�<�~�8{���g�,
"H��Z-[��+*�3\��1���~/�s��K��Z�#qܢ��&�����~����,tO��
�0cبu/�(�U9��Y����Z8���һGBԭ�g�v`��$M 	/Ơ�2�K������N�ևr�ބ�1�ī�,�k6��g�^������c��%x�//EX�{!h��t����;
01��,P�<����.p/|� g�t��q�)���od��em_Y�'�3l?�熍���4�pm&cĘ!N��3G�ێ�����s�j�3�47���~�B`Ts�b,ω��-����s|l-��r���X�غ7:�G!#��n.y�8���)wSj��C�_�*{�1Jʟ��Nn83�sԼzы�ɕ��F��Z^���K��Q}�i�[  �l�$/m��D)�HH�YZ8�}��]~3�=�"
=@�q�����L2e��PF&�cr9q<ҋ��d���-T���O�����)Y��0a�g�ܟs}ρj��`�!&�mX~��u}s�"�M��n��#ꀺ*���}y������s��I�>%J���d�_#�=�a%oV5������>�P(�ph�˙?��K�rVm�/�Q�g�2?�e��gɏ
���xk��f�N~]�����hE��2*:XF))9#��p���bz�3�|�~Z����16���`uLL�_�����}��H��^���L�}��/�!Oo�?�Z���n�����kG�_qW�}�V|��y^]���t��Q֍A ��領>{I�P�c�&�"r��,�R�S�{�=^��?^��q��[fy?���k\���r�|��F�]�ߘ֤S�_z�6�h��5���S�v�qYzM��o�5��}k�noǙ���Y<�C�ƕ����/;�r�T���Զ������\9�9����}nH9^y�O{=à�'e G��|s�iɴ����M��f�_�X���a��m����r!.d��C£a�[x�Pռn���[�b<���L{���Oq�U�:��Lz��F�U�9�$�:�m��#��M���Q���޸Oدm��>n���[j��Q����k�f���6cbZ9�}CU�:�s�vpJ ������s���oƄ+=y���W�%Za��<Z��ڹ�/2Ƒ�K=�^�������gJ�V���A��v�����K�#�ߦP�Pf���p#U��.2�ϛ%n�TsNy�v��~ͯ�w��=�f[�p�<���>S�١s�|	I�&ˡ�P�	�[�\u$5��1߫�;5�������}��;�l� ���S�jGؙEzI���F��2M��s�7�9�/�d�BBr"bƞD�A�Tn�V� �}��t����s�)�
r���K���F�����H��hDov$ټ�,]l��>�9�+۠����z}�n�H�ȋ
��ʈ-j�"���qAl'��%gA0�ϸ���_���K�tt�_;K�*ѣ0�dh�2X�ęs�n#܉|/7�@ =
��
&��G�t^��:������Pa.&s�:F%!]�m;��pc�[G�'&�\�`���J�B�X[ִ�7ϲ�^�H��+}l��U���;\��rg�w2��[<�b�;jo���=ryCg�-���d;�q����)�|V-8hޥ�C�,�XVXH�zG��I�.k�4��{��Cw��IG�篫qK$�RT���oȴ��%X�u�2�BE�#!R���k�J\{@��p�	����(��j�9�|���G����Ifz���V�곾��ϒ:�Z5��n���V�܏]�ֵ�_�a�����lN�f+�d)�����(�o����C�;��Ȭ�0���k�	��_:&�lcH��ly��:�~Cn0�޶H
���\L ǁ���b( vlG-�w��,�������_�<�����m2�;���}�#C�v?���9�K;6od�mH"ÅV_	[��A�|��l��'iD|&mn>S��j޺�����A@��M-ox��v2��߭0���v	���� Z�՜7�dnP�7�|r\
e���f�F���I�>�Ev"Z�$�e��9�O�8^[c@0��0�UU�l򎸟�"����������酕ge�/�Xj�q�N����X=;#�����rP9s��=
��~F�U���q�dd��Ё��o�����v����ԠayRjU�[X,Q�D@�O�Bd�=��l�fF��u#�� 6O)��%���_c+4�-�E>qڋm�������8� <Hd�߼ϕ�Q."q� P�s�pG�	�#̇�wq�x,�Oi0Ϻ��7Bf|ۺ����*Z��+�eQU�";[�=���f;�3���-< �E���p����( Ԋ�E��J�]����ec]�B&�++6D�d@n�p�ĄH�V/����9`m��˕�F������hkk�벽@���<�
ݢ���aT�0.a~���V�"����E��iPnp	�ǭ��beU��+���ddH/��I���?K��N⯢I����DU�eR,*���8(�H�j�

&���~�c���՜��7s-^,3[��6[s7�h�,h�5J�9��
���k�*N�����3�P��)��C��`�nYD������w�CZG��jk3�j�������{Wb�4��`I����B�Vz��i�����5����G�D�t1J���$�f�5w���M|v08:|�����t�7��p�A�R'�h�d�B���(AG	����-��-\�FA�b��j@BԵ	
4�˝�V"x`kB��]��>)��;A���0��A߶DZ��t�@C@i�C�_�*��mmS離��i*��-���qI��NS��Qx�����>�TIB4EC%q
��=r]>&j��Oh<�u)c3V�lb5�S4#:~Q���}�F%���R��u�DQfG�Ǻ�B�<�c��	�1��^|�r�v�X��w�3*��V�����BPN��<fY��=d���U���S�1��t�K��� �Q�l��J����h-%�CWH�~!�*n��v̞��ݶ���MP�ٓ���h�i��]�����Mg�ITÈ1#XX|v���j��lE�r���,L�Y����6���v�g�������D��bK���J\�M3���q�H�~a��Rx߾$�3Z��Pm�slӂ�O x��G#����u���A�L�����F �C 0�*����� �]�.ߋ���E�E�:]e���R���y{�2��Όߓ��x._�z�At�f�|������'��!��/�%4<����-S��A%��冽y�R@�d�rL��5��E��BlR`	�|��5R�^�7��l�1�w)Ӡb}�0���GD�}ng �Ɣnӧi�F�l��H<��j�R d��$R0�?)t�1�=O���7^�╍�2k"��џ<�L�ݿ�Mk.o\�Y[.��jY*������a�M�M2ׅ�$�~!�	���0�Gy����]�br%/�|��^;��(�� &^�<��1��p����Z4�`��F6�T7�k��G#��p"�D QFz��j[�z7�G��n�cpS\� ����&^� ���aM��k�D��v*V�@�mù�("	k���BS���od���q_?��9획����OP�B�I��+rY�(�l�:�����zL�"O3�*����qZ|��u�/f=��`�b��@æ� #q�]k�?a�)~�򶱄�h0j՝gǮ�#vIdShIs,���˗����A�PDz$�~�%�����p�-�C��G�����w~Hbn"+G"$�w���_k ��[d˻�����a`l�����_!�����Gf~0�/g��[���	AT(�jú�(�U�l��g4��ul���+��^y]֑ex5��nLpǐ \"�.���u�RYLA�, T�3.݆��Z�q5(F>(���:�|@��ٵ��}��[���LN���
�g���	hh�ҳ��t(�T�HI�)9Wq�����ק��IP����V��ܡ!!���!:,�1�	�B�zj6�^ ��c���I4��x��$�4���O�k��JG���@ރ���>�K���ӈʅ��B;u��{
/����S2���B/���{��	_n���}�����
�d�T��ٳ��?4�@a���]��*�(������O���T�ȑ��`�HU\=yr��Z�X��an��CdD΂�����4��5�#J�5C����D�48I�]r�n��r�x,�
u �4�w4x��"�X��S��*m4W8- ��$��+����}^�.}���"��l��S�M��pP�N���H��+�B�VbKq��������Ҕ������n�.��R�b��V2@G��=~�a �\-�BA���b0��>��� 1���5����A�����sC1��� �D�;�7_ r?m�4��~����7H}fx
���~��Z���~M��9��.�*�nk�x �5;�&�y��*����+�`�T����K.��oD��x�7$�ut`==á�b��R����t6P��Ǐ�B����q��]��'_k�R^����1Mz��z��Qf)��E"����4��C0C�>�<��yE!���rK`Y*�=�$^����T6�Xɗ;�%�JA[Ԩ�[mH�m��Ph"�-�$ݗ<�pt�)H=)=:�d𨎿N
1��߯ 0�Ej��\�팷q�q����s��p��.�~�b�y`Aa[4�J������"Te�CP�����"�9~���=��g��9Y��B��[&��Π����e�o�����-�3���ǳǾ�h�UE���9�
�ʐis�Z)�#�-h�W�� '��]2D���&���Gƪ %�02sr$��(i�d\�
�1ެ5����(���X���ڟ$���T�li���X
�R ��"�o�l�FrPQ��m>\�MW����l�cn��e6YT����_I��8�����ⴊ�:���)t�tj��"2�J�ۗ�ǃ���������Hl�K+~@΃�Wh}�Wa�<�4 ۿ�ݲ�3i�"�C'*�DT�^i.ܱvۯ���>�0�B ���z����=��:C嗣&�&>��C$iy��>�<#;x�vwե����@�]x��#���<孷���j�x������f� zX�S�aB�&u �z�!�V*�$ UO��b�X�Vf/�l���%�alBF����騜U��gi���>4�kjj��Q~92�ߒ���HT2�e�.�X����# J�s��y�l@�4�. ��4k�&��>hd:� ��6H��e����h&��c�T��b�9��t;#{���#��y^J$n�h���z����J�uȍ_ݠL[k5�e��qH&zn/����A�|�����������<��a>�ջ�l�f�}��py�.l���R���j����_8XW>!?��$��i����s�)Զ�u�+o����6 N	�s���ɀNl����l�jP�K3��Zt�TPnj��g��9G덊@e�(x��[2-�HY�9�Q:�I瘠��:1ǫ]�G��0T1�T�z+��zf�鿻�4��٫8��K�~`�F
F/�0!"g��D�����}�5��Kr���3X��	�2��uv�趆��S9��A��Q��Ȅb�L'l�d���~�]Ҽ�t3�~��O���.�>H���>9�Z�j���l���c��l���؛zq3�O����f��o�cي(+�~��gVB��2�K�)\d~�HHA���|�T�%^
0g`G�Ĵ�C,��B����[d��e��w����w��7���1mh�2��f(���Y��m��xs$����9�lr2��-��!f�!7 l��I����N
D�ٽl�7�K�Φ������oV��� �<�.�*@0�{��i�E�����\K�meߗJ����]��.	������?RPHHIHII�ʯu=D�XMՇ��ݑ���A;a��!�ZG����%Wi*�;/l_֐R԰7 *$OE1O�A� 3�&@M�
{�G4sds�]�a�VE���
������l��� �>�Oh��eyPJ]��]��Q[]�,��o��b��v��<:e�-W�Fɚ]��[�a�Ҹ9[� ֪�=��Oz4#�l�lRX0�K�1� ��z,�4ğr� h�V��� ۏ�"�-��v7)�Y��zRH>`+~�wfO��A��#*_|�7��wbc�I%�"�h^`5Qv�{�б�����8�e}����׸#h�/:����t냆�ҲI(p���k'�&�^-���H��<��}o'��S�t˟tuu-I�ɽ�ɋ�P��@��v<C�b���8�j��d���ː���w�j�4��ٿ�L�I���m0$;W/�1�@
A�V�p>2<,��H+<-�Gl��hM�'�f�)��b��N���#4m���8����B|���K&��t�8�"� 9�L}� =�i����+�b4���\*߫�]̙;������h�ɐic� f���\H���0~#���:��[Da�9�hSq(�Ua1��R����1����M}��@�5g�&� ��m���'<���rn���oR�#��6RZ�룠9�!Sex�p�C�[hwh��UX85'&���'?�����$���:x��vҐ݆�mG��o�H�|E���"��X��~��l�``�@S�����h�X��΀K�$Z��s�X@���U�H��br�����E0/!H �`h�3���a�ێ��O�j(�P��%6O��IE����J�� �0�p�n��u&�Ā���*�}
H��_ł+!�m��݀��*�c�@�+�7�����l��X6˭<�;M��$�n;�e�x�Z��g���ԧ��Il�+�F�m]rh�� 4C@AF����a��6~8
�#`f@�7�)\0���4���<�P �$��X狈^��a��� ;��n�"�l���-�yy��G�dn��� �-)�~�r�x� ^��?ˬ�a�i ��Ѐ���L�138����4�����j�Ρy�l�h^��������	�J��6��Hb��!���`F��i����W�7E(��Rm>��� ���^d9�p(wt䙙~�LGճ�d���	A��ܮ�꽏�����{�;mp�6l�R�1���2��_{e�Jv���(���{ ,�U���!����)�X!��ܚ�(;�~�2!
�����Iyq�E��ݍX�A���C�sw��\T�d����~���9����5�)�l`��90����כMX��[���r����"�#ض̆��r{:����^��z8��Z]�r>��|�
���J��z���ɝ�H���������_�X�x�p���>V�3q�S�WP�T��S�����v����L��f���wu.��V�{�v� a��������g�L���gVi{��,�X����9]K1v�����κ��l,���:��.ju��d��&�Ϟ,2���]!���i�.R�U�i�B;�mFf`�+񽮸ѝ�u��q���Fh�c1N�n�Ϲ|;?���b�i�n}�	���,c����<��O�$��|�5�ި:86. K��I\Q6�yc	��o�r�(hIƅ��A���W�����}}�㥠=.���������m�M�
?���;?^��U�G�~QR�����Ix��	�[���+�_c���8!p�9����y_����cp�j}��p�PU��if������4}�������y\-X~���Q���@�ɝ���+���_j-���#�.R�о�[mkݶ���P����G߉cU�dBǎ�����t~*�_ʨ����o9��M�� �g��r�w���5S�xd�M�����C�zǫ�A��k[��w�H�Fļ�h�Iv2�^�U�+�Ľ����^��00���k�׉)z�F�UI��F�=Ӷ�׍hw�=���\��5dw�v����Q,���r�����;)���� ���2���i[�E{�|;�5^�����9�)�U�-��}&ZS��k�z��樿U^�~�dp�d�r4��u{CJĞ���v��nG����K�����:���@�s�{G7�:���v����ކTW[+�����Qu�[t�I�jG�s>�X�ٮ��8�hEn�~�pGl}Y�_�T<�{�~��\{Y�N�&{�� ����dx���Hq|��w�_�mџW�OZ��%�=y/%�;����W]t:���ӕR�ΰL|�'��P���r#�-F����5u��7Ew{A����˖�� ��yΆ蔲�k�b��}�xû�����Ҏ)��\s�q������ֻ�ޮ}7������:��'Qt�V�7�9WB�O��W��s�.��Km4j����lfD=�MR�6j_��16�-���[�v��7�ٵ&>1U.{��T��AY��u��ߛ�%�h3j+�������'%2��:��X����kk�����KB�2�}s�f���������'k셣k�4q?�8���J�l�%����*4���6��aN���6�P��<wĮ�� *����*7`��$,u~�p�&��=���B��/�;"}򑢵����*=�{�|ԅg#�Ѱ��-���%�$�H<ߓ9!�fd߳.ץ�Y�fd�W�$s{J��AM&	pG>>4W��p��k�DG�l"nsE�8����f�M���3È�' ::����!�zafn!p U.�������f
�=, �+y�e*zW�g zqc4`!O�Gs{��67G����z�&-��r^J���+�$ex݃� 6�_��;�|�}|��wW5p���?�;��+\Q�h��K��L�N�|��滸�5��`!�޾ߴ���d����l�8�V�{����W,�]]��u�����(*	Z�o��NQ�9�/�g��6S�ÌA ;�fM��3$`W��\=XhQ1B��m{�=�:���$z_\i�{k�E-�N�ɣ�����,��:������L����*��E��;׾Q	�� ��(�8(�G<RXI-�S��ߒ�6����4�\��j��|����CL%1�,i��J�sP7	����>�i���R��K����ۻ�M�)�g��p�ܟ$����~�/���z�Fݥ��HV�Cj1@
�]d����V�W�I��l�X�
)�np��\�l�˩��oT�aaV�����	9���Ȣ�~����`9�Ǧ#�M�Ǯ��.BYu����������cH^ �74�g ��eEFwzb��7\R������W �$-��κ�D L���%b��	5���n�&�[Z;)�$1 	��3A".�[?��
s�^;��/�Y�@x�VR�����0;��/CO����1R��
�Sw��8|U?�b��g�O�-!n�p����灒£�?����5��fx��4y�g�Z~��yU��`n���=��x�>��¦�*5M_6�﷿�o�uO8u��OuE5樜>b�94���+�n8c���+R{��|�V~N��j	9~�on��ڃ���ѝ��Jg��(�%����]U��yGc�[9`s^nJ���'	Ԝ��6�t8�Z�ޓN{��6����,*~
�̸�zƛ���P�H.`Dt�vBD��^��DI���S���-O��PVڽ`k���Y��C��Ư#��w��ʮ�u�,�P�jGy��ߏ}��ke�O~�捎�6�5�)�֢����zG���֚�����B�r�"XQ�o��uɅ1fXo��PX]�[��7l��pY��6�I��w�i�z������v��J�%婻oa�E�=]�.�~�G�r�?zJ��4r�H���i�00N���#�,Q#·^n2����6���8 �$B�@�L�}�b�^W��(��}~��dZ���s��Ni"��Od��I����%�8���/O��/糿���?�sK�~w/a�e6��U.�"
���n�ϒ�hh�b�a??�\���h�Q,zG�S��`j���)�~��
Z�y��fѺ+����#ꆸ5�ݤ"������sLWy�������qP'3�T�F䥝����(�4��X�~��l���ğ��t�,�V������]�����W��G�85M�.�F⟠�heU��p��}WUK�?�ե������P�U_[ˌ�v���.b�+n)�n��<�]��?I��$�@�V����uճ�(�?~7��L��uX<�p��7�N3k15Wk�[��Ѿ�k��j}��Z;n�h�?�н��8�e#���+*ԏ���Y��/��N,ե��ȼՈKm�G2KҎ��������3Α��?��SRo x�j&��Y�������1�����\9I������Z����:LPЂ���"�>U���	�*�����O���'�ӛe�y��}�Km���gEX<H�w<n�8c4�eE�H��������M���XZ^�֖���=�3��P�� |��������NI����ZoT�G]��kn�6�t�ܑ�Y�����g7=��^!�늀T��Oq�s�B����$��l��c���/����,R���ѼՓ�]����>��3��(�[a��@܎�/����N	�3�}� -^�h�x~�� �Q	��X�%�/)�D���ao��S����o�y+`p����8��Z�΄]�ُ�؀�:�%���6�.@S7��G��H��.Ȍ���<@�J��e�A�>h�#�'�7�;�ǫ~�<���+Ϭ
_\W�~ݬ����'�~ʓ���l� @dx�uk莑�9=�]�v=sH�����m�ĺ�%�\����4w�Oy����g]xz��48��`�[�nI9��z
,��׮�]{�h��l����o���v�����޿�~�ޘ>�^�Mx��i����W%��ȍ~����p��)���%Ĩda�'rh10-M:6i�� cfA�)%5���>� �y _/ ބ��N�o�1�r�dg�o�|V��5"�ܗ��]�k$y�2Y�Ji>�#��A�.6�H���_�]ND�H�~&����@���@X�����T���c6��fܴ�R����\�)�C�l����z�=��QT�\��V_�x�죵����i�\��.�,�f�ڽ���2��"0����&�Um����T�OdL�S��dmMU�Q19��(�c Y�<����<��p��w;��C������bzV����|6z��Z�0H�AW!E,�8O��Q�F����Qƪ�&,P9��9ƠkA5���rG���W�f�r��y�jp*��~�%��CLP��A����|w�����^��+d�C�~�	?%��d���+e�2�I�����o'VL�U�M��W�?��d�]�{�1K�i��J�~8��sᚳ��s����N����h��{�ㇵ�������{�QA%DDZAJ��K��E��`�!DA��`讁�������{b�O�/��Ď{_�u_�ޏ�E�WD��Rx#v�n~�w�I��)��tR�m�}��xFj�tߴz���,�%.�[�@1>�.4~�-��]�g�uY�d��؁���|BYfB��?�,G��{Kf��d��IG6���(g}����"Sީ�t��eyGz��]]�^�~.[AAM�I)g��@k@zԥD�MQ��L��b���c�D�`_w6�U�f�����9�޹�ܪuW�}���4S�"�L#��J�#!Y���r��;>O:���E�%=��i.k���=m�@�1�ː��:46T�@sQNoma�^�M֔��i=�a,��;h�AY�8��M��@��pM�������C@R�j�>qZ�j�$�i�����<h���1x��L�pM�/���?��K�(�^^��T��r~18��~� ��#�HƵm+��F�: #ؑ��0Q�6�P��)���W)&l�_MT��,�0!`kG��^�������w�����i:��,Y�]���D�(�m���I1f�K���|!��"�e��ȝ�	'�WǵU
�r�ɶCЧ�z����@2d�3���BuV�n�}.����]�1T���8Ʃ&k�>���Ī0I���ًY�l���9���wQ�K˔=��-�x[0�6��#w�����KX���_T�f�S���i��#����_�x���(������O�~e���<������7!S�xSd���B]���B�l;/[A�;oWۨ�t��ݢ�����[ߚ7���9>��24$���G��O=��D"�Yyޛ�2kui��b�׶c��?��Iې��yr&��&uT</ ��"�o����7�}.'�j_W;��H�1ez�E�)fd�E��	�͋�)~@'�ǫ���z�Nļ�!j<��"�@�����۩Ǜ�i<[��_�}�J渗��-+��g�"�Q�vIVWF������C����a����W̢�Z�|�&#�p���X���rb�˚�=Å���e�	��'�Q,L;�[�2�_uE>,����}�=�Lg
6yx$��4�$�5k�A�8�|���]����&�,]�c�u�w>����.�~�ъzM��bi¹[��R���d|×'��(ݽ=��䡯�b�����7N�)~�I�$_<�rW�u��划ĸ8��Tt/w%^��N���A��bs�?}�"�	x`�ř ȍ�W�����&yDh�_��:n�����?����2�`��Rx���-G�S�Ǩ�L@�Ȅ��i���p���S��@��j��Fz���Ț�r�P��;��|�w6ў�r�NxkBN<�Z�NtP���$�jvH>�����~���`<!���ne���ځ����@�����]�:!B�1����!�s�m�Y���r���È���mZ�Z_�p}t�ޛ�f���9��"�Ғ\:�$O��pg�>v����k9/��B���E�k��Ne ��(�`v�E�$wt��f^�]=U�Ć�Q�S��g��F�ٳ�y0��ލ���h��1n�
��N��(E���<��7~$����b���g_O/f�N]q�hH[���M̆�# ���� Ͽ���]��>/���%����EAF_����)e&wa]hI|h��eߛ���gKk�J�mׅ'������ќ�%�PO1��g�@��2�J<m?��F�7��t��I0���kLdr�~U)`s�E� Ѩ�{���jIɉ=edXʓ��.��jq�����Ͽ���xH4�ڨ�1��p�V7FO%\�!�E�̑�1r�3`4/h2��������Um��)�R���ߢM�_�}�S��Ҿ��kbN��[�T�>�-/z����ђ'j��x�Axη_��Ʋ��a�a���^V㔳f$�h`��׍�����q%��jT�L�J[d�t|���*�z6'�db�/(�'���d�d���7�`:q�e�R7޽[�ʲ����Ҧ'��N��#m5"9���0���ߠ�\��KzG���G�Q���F��b��Bun��Rq�J��s1'��3z�(8b2���R�`oX��q��
ὴ�k��Ϳ��?o�a��\�3ct�a��Ez�/�P�(4���5�S�7������]�>�V�T�+�Da*腡��̊=N(��&��8<H���Mdޅk)�n�l|{�������{~�����[���y�X>Y%�����Ԉܯ)�I�\'I<�Cwv♩��BN�����b�ĥ�]A��#Rb�6���[0��n^�
��r���@�)tnӛg?�H�{{��I��/ͺ�`T~�ۖ
\ڮ�-W�|r��,핿c�X�哗~!���nS���ܼ+ho6da^���4�#��n~O����K#���`4%��溧�8�Tm��A7փ*�5yFV
[����Y	i�ya>�ˏ�4]A�������Hp��i0�YE�{��,4�ڗHf����LÈ��;,�� �J}+OQn>�gh��xL��X=���{j�+#��ry�]gՎ�rO���f��BF�|Ԍ4��H�li�e���%�;7�cr*��疝I�W�or&�8A���+Ku$;��7�RO�ao��lr�!	�|�d5�몮]y�ѫ��d�C.���;N�'w��l&�v_��{�K��f�S���/����WI��X�r?!=dM���X�i�.�����I^�.Hg�X�9��rY�+�S��T��g��L�wc��EX�MRV:������lr,�.��M���3N��W��t���T劷�/߾Q`
"�%%��S�u|���{b+���/�dz�6ș����ʓ�
�e�T4�J60ٶ�$0F�#Ll�C�\��^a�,1�'tҖ���Reu��mn��mޟz�M��od�7)�klu�~��_�X��4/�������p�D��u\_z���I�W��DX��HWl��rto�o~e�)�lh�96�$?��F�^@����م8/;�ћ��\�k��r�<�m\f�y���'C�*5;�:��7I)����
qtY^�v�X���<�� 'B�1�V��w�{s�e+�x��+��TK֣�v�e��r,<=�$$$�#�C3W��m����^�����J��UD&}��������Ok񬎑����+�!�dU��Zbo3��������U�Ӡ.�@Tп���?��n�������?Y�n�w�i	��pI�q*uv�*��	�l
M.z�"U,l��c�l�}d���6	Q�#QHv6q��.��Y�daN/]%\�k�F���[��:�$�K�����Fn��Yh�b�F&���.�"޽,q��#DOm7�k)���6��Q+�L�(#��(�Hg\y��VE�H�S��'�?ޫ{Sȁ�I�S�F�n/N
��&�Cf�ɷr�]��a�_,U"�^��Z=��r>�<+z%xr�X�5�0&Ȳ�����p_`��.(��o���
���â?��2D������7�V�/�����_�ܸ)o3k�n0�>���W�8�qB�Ιd� ۆz
��	���[o�T�UK�o,��ׇ�v�������W�,eb���W
9X��%�b�aϞ^�"�(�!/}�c��&��M�7.��|n5�?�F-�E;�b\_�*�蚳�5.���p�=�2ȎR�ݝ������z� zk1-�y?�+�E��a}
EC�M�'�n�+^��3����h��hA��ُ���>6#[UR6�9J��D)�19�<&�kC�� ��ti~m�u
��X>�]:�mۏ*��_$6S�9��?���=�k��N�+~���o���*�53W�ޫ8v��L�P�с@,�����h��jج����
`dq��8:�s;�=D/$的<�*�����JTW�y�V�* �-��1�H��29��M��(@;���� ��4]���7��w;v�,	�9��}��p�*<���p���˛K���89�����u���7��I'_Zjn����ʖ��������$+{h����tBI|Lx�ى�r�W���˔�P��$?!]=���MY�F:泰�2�>� ��Du�M�tb�rr�VnKW��S���,ƕlUفD�GS�;۸�&���������5�5�h[H�^Q���O�fMO�-J-(J�ƽ��P@ (p����ξu�V��~5c��/�ˬ���f����v�*w�ᬩS��=���}���?Y�q	��U֗Wg45�P%�Z����]�p?�����Z�~	���i�y#����(�~�y��K��^ڮ,HB��H�9�|?滹���s~W=�m�$����i��Q�]^5z�c��V�'���r�p�^v�5�z������>��)��|��(o'�wR{�o��8��IИ��I�r���ξG����u��ۼ�4�l�0�+��	��eD��=@���V#8w_��?*��_���7��ųr��0�������>�Ye��WTo��x��1��%�� �(�`�z��/sI�D�o�V`U��3N��쌉�u���5���ŹĄ�?�BJ��~���ؕњ�;2��Ns<�Z�y�i���r�_�)r�~��n2�2�SC6�$җ�b�����t������(�ו��0(y�k����덶Z�H�
��'�K~(!��]��-�h�(�I|<�㓟��H�$���{y��j�����-CȄp���[���Ȃ��"�>����SX�\�����N*Q�ȴ����b���[؞�����]c;��I@O�����0�̭�K���Z��&rٍ|�JXc�L���-�<��t���L��������8Zۤ0�y�~��"�Ef�ۼ�xc��r��<�̬�ץ���q-�(��\nc���d��I͟z�4 �8C��篸tH��/�AP>�ii��0�I�SWEw�������j���(	M|��+���})Mr�\\�\q�}��ȝ���d:�{h�V�.�h�cx�#\��b#����|�+zCB�[+Ȼ�>���W�G�u�LT��)��_A��@�|es�n/�cut�:'|���Ǎɺ8�~@���zP�j��ρ����׼�O�b�R�c�����Y����	�o%<{�|&Mwo�B��|�g.d���(6 �9��i�!h;e��KbM�������"�ک>-?����t���Y-�=QQ�4����iN��7�(b P�s��ݺ�����fe٪��h����H��Q��ǎo5�6��^�&�)�� �e*��.���6��OҨ]���0��#b\� �1���*�?̂�1�oS��ϫ�?RB:�.�k��yR��[�s����=��7ys��rj�L<풐6u����zn�>)�SlQ���_�[:����uq����������_�,���eH�TB���.!|3~�������e�SB<h�`?��*X�7��3xD~;{�<�M��M�0�4����/ �qdޟ�ؕ��W:�'��ZIAϙ���hh�����2�"?n/�!#�������Ȅ���>�ގ =�- X�է#u��_EJ���c^�r��wA�	�$ê�>��J2�.)��L������`����l8].�֪��[���7��W�����k!1��v�u���X�=�{_'�X�뷓-C��N����g��
�U6?!�Z��3x�&)��^'�����xFv :�/E]��_k�\�������S��>�9aF`2�Q&i���_�-�o��mR1KS�5Сٝ�	�|����lO����r��Xu���>j;}�����G���tBE��	�hzP�7�@�i����]I�]K��F��̭9�W7��]��3h����}��mKww����SE���Q�w�/ۉqv�\K�b8��è�52��=� �|������Ƹn�w/���hD���	��x	}w$��MG�vko�Ę2m��7L�t���ӿ�Lս;�t�RK�&Å�t	�I_�ʹ�V�i
��������V��x�x�jR�f!��~��C���̇�q��0'�������a+ϳ��})p/���U@
ܽ���<�
b{ �V��-ZB'Y!�w8�v���A"�p�T� �D�w5�+D��g�[��۽�Phཅ`u�Ut���T�'ٯ���- $�K�7)���8B?HĦTﺎ+�
����7��Ueܭ�?$���p���~��r[�W7+m����`�ω���@��4��;�ܚ��8�1�ʅ"��v��^.�/1YAA:�6��|:���

�~������Ns�S��gϺ#`"%�/�� E��r"�v&^��?~�c�_8��,�J�>%��.�q�����Ϝ��]�� Y�-7��^���Zz.WZzl	��ȱ�\�b��è�uC���s&�6�� ��=|�R������@���
r0�lu��IF�?=fb�R�� � WzH��JV:7�E��q�W�&�Rv"v;��;�3����Y^��<�.��(��@�䂇�F]�J����f�?@w��(N���k��2r�_�� +��,�С.�q~о~���V���fN�6�����NG�'ci����VR-`㸫���te�Wg"upɣ��Ke7�ؽ�q"W�,p����ʽ����b}�k�H� ��C����\�����wo�Qf+4��"�-���K;5��tq���c�J�|�l�Q���Y����t*I-H���zO�l+K��h�UB�c���ճg���\<�r�rS��}�H��n	n�U��~����b.g.��je�B�F2b�?��%�n�\�tV��UZ�@tP�Rr�ټ�!1 !b&r���Aů�>;�ܘO=�'�_<��p1�������ݐ!;ܪ�vn��80h�q�m7�����>��!lW��kUk�<̣�b,/v���`��S[�:G+��P���F'w��c <Z.X�f6�`1!wْ��Td�;��O۠}Wp�EC�~U��ݲ��UE��z��7��/�?M�M��El���C����e�� �� �|8��!f\��ʇ�J��aѷ+?����M� ���1U��EXCsপ�����;�e�Q&)}��m>�w>2�q�����C_�P-�5Ir�]�o�I��[�!���!y�ڵ=_iқÛ��w�Ol�VI\��[���&��C]Z�;��=������^С,�à*A��>`�?
����Ʈֱo��^�+�.D]L��ȔM��C�*@���G+�즶�ǒ_�.�O��{}���u)������Y{��(j�c?���u���c�����S1���^���W�ٞC�ղJ"^�6����[�����J�2��z)}`�j�y`a��4!�ck�6�b�]�x�"+{-A��zNr�"�\`2�}u����Z���t�\��k����i������2\����֏.��	�����r���������|��}�b��8xl}��u�
YNԪ��_B7�(<�-��;�^Oc��^�������O!��<uD�C������8��hB�``�R?�Ҭ(@���q�}MHh}�W�δ/띜o�u�U�+I#�� ��>rR#'��#G?q��<G���Kt�ޖգ��8U�����&��^.�C7����H�PT�*����7m�M��X�a��x{�����w��o�IFHl��t;���qd�]
C>-Rg�.ebe;��D�o+N-/OE�m����m�Ȃg''�3��v,��0Q�U%��6���c(lb)�5�ϬXBF	�.Wk��C�!���*A�j��č|P�]=-���^+:�NK�T�#�]�'���q{�d�L� ���VN �����>=��*pc���Dw�o��	��0o#�X��<j��(�A��B����U$0C9F'���ǝ���u�jO�N/���rYyNɑ-\����Z�d
;��V�6^דv������=!�ǝUȔRW._{��t�C�ֵ�/�z����#������Z���{�.���<M��*|��K|Z�ՊƝzI�B�<k`I`���wU�7Cu#3�%P~��@�XZ8"�M&��f:v���7�Τ�;m�������!�u������]2G�I�g���+���E�+j��t$��{*���=ۮ^����@ł`��Y��,�s�@���}�B�� .���������v�nB��5X��Ωg�9��*Gi�{�9fd�zt0[��x�`���ê������ȫ[�X����-�Rv$�Θ
�����_�H0� Y�r�_���X�D��ݻ�Ϟ���(k��Ctө��.�)V��3q�uEʢ�f��y����K�+>����]���SQaR��KQ�t�ʇˍfe)�T}u�]�r���`l�ٕ�����Ӿ��^��ʗ~���㮝a���c��z�xX�,_n�[���ss������A*]���8�x�m����7V�ը���?].�3GBbJ&'��
�MQo�Hh���8�}-�b�n�O3�ʙ
�4�>�G�̀m��g
�.��H�):=)5�c�$L�����j�tS�f�R!P���#w9U��zNlU�V��&�ʖ�/ŧN49�����E��+��;R���nE9f�����H������:�"�5�1M�x��Ѣ�6N�Pf��ߚ0�V\����p;���"ʀz���m�1����_���Y�MY-��{d�H���x2�v�n�m�4�X��s�������-W��n���9e��|�������.T�k�;�O,�[������o��k��z:�?{�m��YXR���<��K�x]�e��eɛ��s��r�u,:̮��)�'#�E��^��J�aųgTd �`�^ǻ���Z����D�y�`��sz�ۣ���g���`�V�"��Gz��ꍼ��̃
a�!����AV�Do�-�j���RPǱ��}���5ŴiJ8X�5t
E��&��t����]�R J&��eka���.���.e,r��X�2RօҴ� �E1)%�+*{�����:��0F��%r2��-	з9�7`��A���6^���f�-��p�$x���:�*�w>Yb��b��"�4J!��30{���L$GTF7\�e�JE��z}g�A,�O��L�f&Vd��s7���/����c�Ў�Ȇ0R���:�2P�y�����7�Z�&�j����
��������i��S�`_%I
xRC����hb�l����~^~N(!�\�|��ߡ1��×��A�^H�>
Q�?
�5ղ�Y����/ 3|�8�
MQj
�?�wS1Ў6��Nme�G�҅]=+�r�.}�d�CE�bQ��������0���/��S�o�񥚡�1R����?cP\"��79Tc���b)�M�k���ٳ#g`�q5�8D{�(��S���Gps(kDF��]U��C6�9�+�&+�ψ�s�k��c��0G`r�U�=D�ִD�^�n'��-\"��?5��>\��0_��N���U�ږ�ls���E��+�K�~/��Ŗ.��O!Ҟ؎snc��K/�]� ώ쿾L ��p>�Y7]�����#�q�f��O��	Ӓ�hJz�e� fW`��*�� ��,����ʟ�D_
^# ����Q�_�m�/�v]�����X�82�Q��~�f�2W�'��^@����������ޜ{u`�:.��i�z6��L��
�w�,��U��!*'��%,����]�\�{>ԋ|w�}�Bޟ�=���9. �ݝ�-Slo�+�3�^V�9B,x���x����d���5z_-K{��lt�	#J#O�ٗ�����e�~4��v9�,B�:k�IW�6����r��k�voل�*A[B^�b��R��v��e�o.����N�QV�B�,T��LF�+��u7S�QU�BnS��ߏ���nɅ4{۔
�=Tƭ+�~u*')�W���ͻ�?�m׉kb��`���+j�yŬ=���r�[���3,/y�+q����F=���T��J���3#!v��(K�m $��If�8���L�E�([J����[+S�����
��8f��޾|��-���_����a�ź�({:�(q��D��h7?)��ЬtR�9��V/�%vcZ8p���Jf�r�O�D��q���m���3���)��;�_��P�U�`鵰�u��n��l�����7�����zUTR�%�?kB&#�gݷ� $;����xX+W�ʗ�AO��//���Xߕ���p���'A��]M�	���~���q���z+���{#^��h�ī�g�����Ɂ;͗�%�� �"*�.S.kXki���Z�1��*w���-ъ鬌��P7��"�U�,p;����h�<-%
j�].4h�<�Qh��- ��SN�T0��Ȥ2csOӴ��V��_�E�z��6S�SH%�>�&�� ^h�ѻOx���ֹ�|�&O����M�`���Ų�Y���߯�w��C�}�be�w�yz�E��"atP!`L��P���Oυ=���~������c���@���R���o�Y	������r���X#�6w/n���D��pL�v��f�8n��I+�fh���9�㉦�鋯�x3we�/���~��\kR�@�<��$�|���g_�+h�ˢֆ���9�g�?�IXQ�R��������1�%������!*�t��_޴�L��}�(�l��'%X���;sBx#�ޝ�^豬�'3��T��/(\���P�K~T-��Y���y������[�X�
��]��߸إk�g�V%�����S��^1X%��W�}��<��M�"B�p�1�s���i�x�h���O0}�c1��{���b���@��Ǳ���6���E\`0d�\)mqF��#�f�������4�����ZǲИX {j��p�@���ecY*덾\�}��<�T����g���[����9aa�y\J��U���(�v�W/k�,lx0�.?�%��|Ų���gMZq����e���0�$$��2e�8"�;"�,+�-�P
������a}{��C8%nr?Z���� JKN�S}h���p0S�������������{�)B�^����HEр�ۗ*f��u_�V}@��x識	�� E3n(����Y|����nj��!l�Q1/Z�z�4~+�|l���4˓��n�qKe�(� �Vd��;��S_���iM�"���v{��=ܬx�:b�g���by�I.�X�n"_��Y��)��?�`�Ih8ǼN�?�#l��i+]�,�,�~�9=���)���b�w����N�?��K�����M��uO�L+�߇���Q�g�:)�(؏�+�>��/1m#)J�t-����iTe�˜:�eӉ����/��Aƹ5��ùF��}�Ug7Q3�z�+ݿ�}1�8�<O^��C[�w�je9��A�y<Z#I�Wr<pTe��B���i҂�ʵ�"�UӖjyZ9���yZʄ������gh1{��{aO��R<ER�c�۶�~�:�����2`+�}����]��HG�Y���ݩu���}Y}&IO��*+{�޸�UbX��x6D�V�ez��"�-�$U��u�0l���l�̛u8���)r�Zس��"j�E� �a�O-����q>�T9�w�>?��@����LL�q���%2��n?��E�FF�a�͋�[�VE@����O�'w0X��KP�0���I�1ο���G����z�I_aծ�����"��2V���g	<K�#þ���޻�|<�ỏ��}�"FV*|�]WT�V�����t=�d+A�O�i�:���$�rƪ��H�=8��h
�����teV�j��pE��fz\�Խ�n��3/0�w�J"��غW4��~�B�eӊ���f"
�����V��p��Ɛ���H�B�#�P��[��>7�����t��x��m;��ن2�ޖ� u/��KBp�)P��,��B{A��5��醑�~��ݛ�oͤ2~$�˸����W2����-��9�cRGö�����@�Zy�~����������'�Ӧd6_#3��ϗ�^o��	Y��=o[�ެ��q�;b��tQ�_��Ɖ}�+��DP���U��	���^M��PСZ2<�k[)��؅'�Y�G�1m�	�y��q*�_zu�=E�N���o���A_\P�1��3e)���=��N�^�.��r>(){~w����`k���ȮJ�YxJjWR�i.���I�f���f��'��VwYs�:ShT]c�;?W��g������������x���`����O��U"v>��`��wr�S�&r �L(��T��f)�o�}��޻5s��/,X|�Yi�(x3�+�JFfωA��S"�}�;r%�g�?]�Hq�Al�hĤ����tjv�q|�P�{�g7/�Ko�,�<e-t{��{$�y��5�����틳�%�YԎ����=mc�ޢ8�#I&�"��?K5�E}dB7<W��C�*����Z�8[��v�3nV�B,���&�Ϥ^�s���ik��*�H��ў���L���+��|#�e`��k$}�}�Ӭ��ìŶ�$J�?r�}iɅ�*��5���������3���_ƈN�\J�]�f�ef�V�P˭��G��`nE�~%DmQ��P8r����ݿO�����$=Z�o�N�MҢ�Q��s�
��^��V��3�_��~NIs�1*�zj>��jى7�W7!�ui�ݘm(�|2����� B�i�[��s��m=����t:F�߫B��⛤��c��L��T3T�ϫ����R�v)m���?���� Ga��f��H׾��ʭ�)��rk�)J�^o�f��:�F�n�	�H���Ӗ�����ػ�Z6�,la_b�D!��ɑ�5Ы��4o��jHGL�*O�0�����S]������>�~��J��+��"��w�Bg���WS-R�Q�0;gY
�P�O�ܻ�Iyz�ZD�z�aQ�����2k֮(��H�=$������Y��p��@�*���/�ػ�v����"{ƾlj�P0������x0iD� ��e*JW�� ���*eZ������ �v��74�ʟ�Q����N��F��g��p���9�<�ߤ��a�ؙ��Q�!���d������C��CC�$ۼ<cb��V%w��y��yK����u��)�Fuǅ ��O�N�n鿅�r��J$��y�Rՙ/���w$]�	���T�%���Q�߂3�+��s����Sz7]���0ePJ��7ir�0a^�Z�{�!�tE`N�5�+���z�@}�I
����5Ǐ�RW�������V7M�����=�Nh-�dİ�_�(N�Z�E}%|L;�
�h��g
�u�GDV��y@�P�v"�7O��9�~0Q�J���N�h�ӴM�B�8��ۖKU2l�~�n?����\xդ"@h
ކ+D����Xh����[.�=��W�7���r��|#��ja
���6������Y=,��4���;i�?�<�w�\��"Mr�s9�Si,"���v��{�M��Il�\o�S�!�N@z��� �V#���/����qj�d�B7�=n�+���극@7t���������;9	���$���(���M���a%�ۨ��Fs�5}���b��4p@8�5 �����귫І���_b�ث}Pm1���]	�0)︪H��׆��?i�D#�Ǘ�
Q��Y0h<�y��Y�)�SQ^` �����-�Gz��pʺ~�$��6Sw�l���1$ +��zE�eN��b�5��mjA3��f[BL�Kw�F7�*jU ����[ډ0U�-�"0�n�B'�ƣf���=�N	́�Y����D�I1�������:������nN��IZl��N
�?�>��Td)� ��/�*;�"��ͫciA��SlՀ����ی��U�*����*MdM�h�� ����7jh��]S���=�ws��+,�3���/�H�N���&��p��p���ti���
��¿|8���f���@�0���>N�
��O��JC�����8�G#fT~��*�	�C�4?�� m�A;�[�)�_F0n�h�!AT�m^��` �t���r'c��I-��2���?~W�jOi��l+ G���J�ݙ�la�m����p�Aİ��j14{�����,͒`�5�~n"���_��i�����1�,J
��6kp��k�_a|O��S7(�N��h�	��BW�������3�z�L;���q�hq1��)�Т��@ZQ�����Y��0��W��ldG�D�A|��5G�]F6Z�?�f�o��t��2c��>U5��>����_��9�-���%)i+�X�OG�O�Z�P��D'��T"��g�����TxM�b8���٨�*��F�<y�hl�.�-�#�9�J����w���_E|III�}�ity���2��T"rJJe---�����/>8��dvS��"-�(�1�iVI����k54��uQ���)Z�s�5���
�;����l��O�����B�0�.�
�z"�0<�Dl�p������y��F�]�wп�����x�Ȓ�4��d��5��q����P��8���`���0�b\Rol���=?+a���X҅ �u(�F?���8�����_
��bV��j���C�9�]E��{j�8�r�q8���GԴ�������W��;���2f:����;��h��ќ����;UQ��<^�����y���4V��#w�!ײ��2��8�,�����G�T۸;)[���	��ꨈ��ƶG�?*"B�2����֢'�Ջ��v�a����Ш3�Z��|�*��������x���S�V���&Ԋɢ�K�����+��F�bX
1�cc:~P�Ѥ�o_�l�v�&d_����^��^��E��PWJ���+�C��Ȑ�!���1����ii����)��B����Y��ֶ����_d0��B�F�0)֘�J�_�5�9�)�
������`p��7�t.��{{U.\ �p�f����H��U�(��G�����*��D)]Y�sz�B��6��[�w~>��ŋ��W�����yP�1��P����+��i�9�Jî���n�8��{.4E��P�ɷ-��>x\`o��j��~��=�N�� B>&8��"@�J~���_�=�I�2-_nn���V�R��Q�`|�x3�eg{�o�"g`p�3��,O�cU�qS��a&�(��P�D^����^��~�ҫ3�L�0���ٙjM�����R��^�I�|��blwW^���������/�x+�\>�z[̵��!��i;���C��Z�B�$��ح>'ҕ2�Mb�k�c�ga��ԙO���5����+X��D�m��}�h��`�Ì�f�M8[a[娠8/
��)�@���q��&��L(��q��(����maj�/=g��V�����Ԣ�s��^���Ȍ��S����_#"Z��#�AĮ� ������?�~}-+h�ͬ��{Tm��,�8[-$$�z��o����в�c�A��!׸}�5fuC�T���O����m��33<��LN�N�s��=��1�� ��#�������p�Y�߳��1�@u��?�d�N���ER�d�睡��s����E�]ǽ7;��ݼ"�/84�����Ν���Ȁ��L.�ɋ�Q��n14Q�v􉍻���ލ+�i�����FY�y�7������w�{�'��ee�g"Us�֚�����[��B�Y_��K���-�p}��]���JIg]��%<��o̊R;gM���4�^*]��s��i���]����W7�p������h�a��j��=s	Q�шg��ޫ�9T�,��b���8}�[T/��$i|T���VIi	��k|w���Z#�M�&Y*���boo$6J:���;7??2""��˩fܑ?I�a:F!;����ffV�+�L��J`}v���]~���!T��]9�T�	ɢRfFƋ���222&\��Ŵe66>�׫�l�lni�`+G�^��f��i�fuS��cbf��eP�(���������ˡq���9�ȱ�Rq˗�H1��o>�����;+��(�x��"�˃[�𸘘�����TTQ����9�rv�k����=7~1nw��2-�t�f�Д����V9����{e�{ص����h�U�2���bhi�i�X�SpgmQ�m�^AᶒV�%+����ohߡ�@��h���z-�3����O�4%'|�'�{c	�$�!��%��-��.��jVP2]y�o���z���@|Lɻ��X�{ff&q3�*�'�J��X���)�U،"�R�Z����������!��T���d�9r� ���7�����(�H�(UQ���g����v]�qq9�B�����eB�-��y���Ř�_r�/�<9�Ⱦf���z�5�����l����/ �ٳ`��@N�q�q���y�{{.y��9 ߽,����Y�V&�_!:�C���x���t%�Ɔ�L�O��fr��ӭQ;�=�noo��`_�{�����$~�+��"(��5�����W�%�����kS�D����۸a�U@E7�����Ł�+;8S{-{t�Q�Q��ji�|)����P4>�i�?��#�z\� ���d���gfeU��K���,��Cxt���~�vj��IQ�kjh�KAЛ���a�gw�b�V��A�
X0��
S�A�sǰz˃ѡcZ��c
�wl*
�E,rd?T�M�Ё()y���1Y�'W��o�f�T��9�����働t^bb�
/�����
����ڕ��^-� R�4����"$��v,@������x���Y�������Ƈ���Kf��K訠?�`�qe2a(����uQ��4-���W��~��������Cu�o�4*6����,���"��J����-<��Ty�p�r�+墬������BL�/W�*�K1
���=�<�?2�#ޫ�l+Y��t���>{D�/6��%ך
��zV�(?�t��#e�!�B�u�L�5h!�3$�l[�{h]� sM�$el#w��m������4Z���Z����T�0} Y�.��qk������ }��	~P�L1�<AI�uwafc����J?8�P!�=tH�Z'��MC���TUY��>�J����\�2Īƨ��D�	h�_�E~H�
z��ݯ_��dq7T�Օg�>�^@B�룅����?P�ػ�� �����K�?��&��0pY��a@u���,����{�/��Z/�B��>L�mֵ��v�]�.����984����V�B4#�m6�i*�ÔO�p���%�����(Z��$%巶���E��v\������%};I������Dj&}^ ෶X'��+W���vě�<��(����S���L��~��{��1�ˮ�e��W<����dA�*��vrDC�
7|~�� �%�ٽg�_��޷wM�?���/]}u\T]-"�tw�4�H
�)CI*�]"JI�P"%  ��"�tww��w��}����7p�9{?�zֳ�>w��z�u�?g�h�mk~���d�H"Gr�T�?S�YPk�uZ���&����X#Z�av�ve���"����Xw��d�^�:�uu�t��k>̄��
�U��%g�����v_
����]p !f��ى����2��_�?���\��|x.�S�(4=]�C���=���>�%<�
�U(��G?:݁)m*7������vz����|��Eod����2�iXe�#��Zq{ϸ*ٽHHmS�J���N-p�����ЌmM��w:�<��xRE<�|N��j�/�%������U`��*��C(mPߑ_�=���nҶ�����Z�_�!ۄ�/}�"�S	D1	���0��-�B�l�}�at��;�5�J���T�2����QfK�w�C�r��?��}p��g�%�:n��o���h>}���ͽ�X2�Ϛ�j--Mz���f���7�~���r��=��I�583	�Δy�Ejzmgn��Ћ,����|<���Ζp܁��Щ������R�|O��n�f��&�N��n΄k�l�aj�'6h��A��4>"�J�%"#���S�A,r�7��/鴺-y\�''�w�oT��~��E���޾ɼ<�_�?W���!*����/O��%C97y��7|���K����k�~L�҅(e�8m��i���M����r��-�[Ai�$6��k�?]W+M��L���8�/�så=��n}����,u����|��W����E����p�W�i��??Q�/�T6#(��h�ْ�R�JG�;-�����5\�e��ؚHJ���}�7�>V8��!)NlDa�9���3C:�ή�>�/�� � r�@���$�&l�G�ՙTooo�p�ZoW�:C�m��i{�HL�k iw��^b�1o�c�Z
�?��x���92��=U���x����c���P�l�V�tdA��ȝ�$��r�{Mjx����6IQ9�WuurR��~��>������}�S
��`t���!�Hp���A���X��6a���d��H�7�Y�
���$b��y+�����j��D���)��+YLo�Y)!��g����D2w����Q�BF[����/V������t���VO�f��#"���}����8A�T��g�U����#.m�郱�>��@���57��j���Wlͭ�.�6��k�j��ք���o�b�P�Dغi��_�����뀋��J�`�
��*4�N��ъ�:`;o.3R��{�6�Fe���lw�Σ=)�H��1q�yW,���
[�X蠺�+����N���xW�b*��y���h��z�pi����ﺝ�AI�ǳͳԴB'����Mn���n��fx�2U��F�d��I_���Zhq�����*:�#Q4���.パ1�ݭѐ�LQ��)ܜJ���]_�5T��@ 4e�ld	�{���@�?�}I�ؘ��G8ˀ��R������_�� ©���f����h�4�ݓm�����rt���>F�)g�^ (A�BSx �Z��1'��?���ĲM�f��<��VDP�����9��G���?�%)k��r�{�g�(�x�ZS�pKĂ��sC���_�X`�C���ۜ_8��P{���mx�Z&�"�{_�O��5TM����\�`�
�8z^�W��x�0�����l+vrr������b<5�It۪������.��;�}��Z��v�o�\�e���Y[�~+��AXDt~|��fBt�8P�D�6ik�8��<�v�K Vq��T�^�9�z�V��|L��{���d�g�'̿�KtYQ�l��J*�a���ޮ� a��8E�^�B��3 @�� �	�����;L���G��c������gi(���MX�������AT�56�F?qX�z���A��<��%`�3B-y�ż�Q������j��:L���擇:��9�~��z�}�h�ZU���eL=U�{���.��Ff�f��gv���9�6��e:���foD\����CB��f|�N���*���=(O�!�~�>e�c��xQgsp�-Qٓ+,��ǳ|(&�OQR�O��G�ύ���r�q���9)))�' �ń������Y�=��'�:�APf�MBm�P:f���dS*>���6��嶯#��{&��l�L��D�啕� %�+���>�m�:��� ����Ὁ�Y���2s��������VM��Bv�;��Х��"%eeK�7��BAGB�5�	�f..�����L�Ԓ�Nu��u�^�4��gW�������������P̜޲!��Tz�}�ob��+��u�,��9�����:�}dF���g0aL�i��%֬X�ٟ�o�<Bղ��
�����I@F�y^fK�H�, )�V��Pqھ��a�V����-q�Q3�W�m��r)��%=�����#7\K +��94-� !�Jfhm��V4K�����4����'<��C:�m
���B4�J��X]��IJ��/U牚;�kc�d �̒r��X���Ub��̍�i�e�����*�'������F7L��&!��+.�p�yi�= ;$uSY�y�G�*=;j�b���$����2�(�́(�ql�)�����z����L@ 1�ݛ���)G_�����`��~2,�~�S��r��������mB�e�fl�|���Y��MW������fNŌ�2����V��sC��Ĝ��~\1bI�y���C��\��)�"Z%b�F��;oWc�g��#���t*�,�͕D:�H����G�yĮD��W�A�`&ϨO�z��#S�#�������\����W�� �lw����us�_�g����H��i23���9�П���!F�V޿�^��Ʈ����{/�Im��{ҹ�Cs��a�Gv��mZl�7�c5��3Ep�ZdogA��m!����ek�#*B��6|V����Nc��;�ĝ:A�+Zs�Y��p�Ą��	�<`��bdddM[e����m�>��94��T�U�z1��������_�G��x>{~Hʥ��WJ}�;`@iy����~���Ӣ�d����w~����o��X���,p�X���z�IAX���p�痣�?|/ҁq���d��������(��TL�[Ș�`i�6��u��ׇ�V���pݸR�4,��&���a�H!n��ͧp;
�>��2�*��׌

�4�Y�fJ֜�C#_v��Ơ��T�� Q!щm���î�m�*�U��J�-Xs+X��W��ٔ�=�T�4d�Gވ�k�P�Dޒ����(�Gv�=$*Q��tnr?��y�L���dɭ��v��]���k��s��x���׌��l��\C�^�	B��!��d`KPP�N� tXNe�[��M��������}�S�>�|1R�dlt4��w�ߗ�I�ϩp~*{o���Q:�<}|ȳn ��g!c�U}3ө¦&����P;f�ϳ�Hv��6�����A�`�2�3s����^FO�l��}E �6L�~傇������K�~�Sz���1M9$���8� y4��k��Bww���o���ȉ���?�U �[��t��G���e]�2#p�x����S�m<!�	��� �4��'tE�����kmV��;��Q�u`ya3ܝǵY����^�ٱg�lOT��/h/|�<�%��%x1�EQ��N�"a���YU�k͟lt���<��y�`+�c�ː��T�k�����|���USe������	]z�$>4�hfI���"	�W;�"�_����	��Q�j�cD5��������CQ����:b[�r6��r��M�1pw�!���l�a�����[����<�i�� ?V���������[(b8��f]�^�w-���&���Z����3|u��]�WT�����ʈf"%�W9�.t�\i��Ũ��y����oN֗��n�~X_���|ck�������h	�KZ�ռ�n��166P���r�+e9HZ�������:���ubf��?}�MO��3�z#��ж�	%����������
Њ�����e��?��5�O���6��|����#��Xr��EMC���W�7P��5���{"BCS����?)qʮ�$����Z\��@M�@-�����{vE3��gf�gϚ��/��pj*m��\o��K��e�D��i�'�����v��_(;�Ó�׏� ���-T��wQ������>  ]��8���2��nK���Z#Q }�(r��%��rJ��)��|�V�}��	��ѥ��ez;�mS����ώ��w{_�)�7n"����2���j5�sIh��ɯ�|�P�ܕvv�+Y��	���^�����a��Ә�ز<���g�x��SP���́�w4���c��sIa�ج�� -~��*�c�G�Â�Bo����{\&l�ؖ�੝�������V�����]͈�����'n��D��	�ͱ_�""��`���D,�1yr���*>Ni��l�Bڎ�D!�T��05��5�k5/,�Q,����6��D�S@����Q�K\n�p7wq�?dkFpD��ar��4Bd.�P	u������HL��<�T_߀�y&�͑4.�˟�-���ߙ<7ܖL`�滢���Ox��J?xV�HH ;п)è`��{���w��4�+Ft�4(D]����V�wVj��*  ����Ն�'��a-��yԛ�[�#a;;;��� mW	/'��:�� �Ŝk�j(�����d1=:�d�ܷ�[�03$�f�j&��C���3���8^�ޞ�8��ެ���`v\�UM���卽ۓ���pD�~l��g�su瀞4P_W��::fJ(-'�E�F�A�]�/�)����=�������ӝ)<�77�5���iH"u�?�4/8�SΝcd^��� ��uA�q�|s<պ�-��j]dx��ٳ��Uk|���5��d��mҰ�����>0�
�P(l���eb��٬�2���`>a�Ƃ�6qp��R�|T�VHt9���?\gMg���g@�kS�}��|p�G*N.uX�I�H�����Bwq���Kt�a��s^*��*�2
q�Iq)��j���N�$�켼�u�����j��ݽ���=�e����?�~�\b����iļ_%Y���{�y����=A�@dd�s������޴cM�c�h/��H}}}�ggc�������]�����r}����?ha�ꝡq���] ^��a��ެ������5P�ΰC�`�'�@U	t��X�7D��D�Z���~��.fNT"<ѓ�!�@�s���UW}��[9g)�uǺ�r22�����C��C=�zEv��ʽѥN�f���2j��L�� ��o}��g&wu��ֲ�Jo�d�=<�<	e�|)v��ZD�yD{�9"m�
#+��\�r�ϸ�w�
Et����1S6ZT���ڣ����͓�4��DG�R�z*�	D�m�=S�p�%�L3�~��Z�9���)n�< �*�[�T�)�[!����l�ht�>�H����rd�y�&���>A�ޒ�X$@�@%w�zAK�%�h�a���������s4�ڜnh}y	i���/����G��^�]��X��/����2�KV}��8-���Y�RlkYsӪ;2��<����L���Mq�ڿ?������|��t=yX�ˣ�L�7��]&۬�5�Y��5Ȗ����ܸc�ͤ�.����2%$�P�Vi�)f!m�ޚ��~M3�{�1-��ά5�#�]r^#��������D��`�J�X�y�N���A���آVc���qR��8
��c:�Z�P��i������H�9P���>�w�U�Z��_~�}�ts��\DWRj��n�����^2�2���*����4g;��GUp�zw�ߙ1m��}=��ĸx \z=Ǣ������c{ȟާJ�׆���E�*��@C�	����$P/��Bk٤��nkL�4�x��z��q��_������GP< DJ���i#n�i�
����k9���襳?�6�y �"��ōԦ����YN�h%��#�������0�^�_BS�\k�m�6im�("CaҠaa+�,"��	�2�T�,�BS�0�kg�c�
W\$蓙0-��?���;Wnޛ�9}�i��3�'r��uQw����"�\��d4���(�t�D�X݀� ���$9Z,@��&a�0��Hqcr�wE��1@����\�����%j�%b�S���`��%S$-�
���nc��F�}�ހ�ڢ�7h�H'���TY 0�I��N��0ǩ�yq���Ah^��R�5��*�^�:W�IN4,T���!1��}��Lz������E
��
C�R�L��@a������3�³��Z���b[�sO �(i����Bomd���C����9�9e��C��8�k!�W�]̶���K����H����)���ې��BxcU��l���Z\E����
���Mx
s��<b�(�'Q���:�O�c�S�_vH�3;�Q�jA.م�czc>�ﺳx�G�S��V�eAM;eSkQճ���N�"�0U��6ʬ����t�RGE���n�@���8���d�k�eZ"3�����ŝ�{Pf�z#7*��T]�Rf5���
�N�Yd�TzuX��
V�y8�F�.��w�dК��{dkHttt�����j���݀�b�'XX�s1�d�����0��54�It���TהԪ�	��f���g���S�R�ܣ�,�i��+i\����I���ճt�EPÅ?u'���*���ʖ����u�v��ߺL�i�Ԅ�O��ќr��gN�ecv�*�
n$���xR�Y�dr�>�_�"���d�\WMT�J,���i��|��K�·h�Y�c�w��z�	-�z��wM����ch� �k=�g��~"/V$�=��/N;P�E��|�R��tG,�N�@U�X��u{#_��E%�5:sQ���6+].��cU�
vA� �a7>fm���n��~�B����]ה.�!�y��w��w"fMC@��Z|��M�1��޲)�T�����H�1���Oi�g����r*�6��'�O�M�Jw]&�~,��˿h�zΥ�mE�Cz"�B$��������Mn�"��?Mi�â=c�J�fҬ_�n*�p���� `|�jNX��Gv{�摙$q-w����h�[����f��2\L�q�]!%��r1�:�U%� 밧����ˤ(͜P�������w
��s�dz��zf���O�����4VKq3�b-V�N��hߣ,�B�UH,��6i�>`��ט�sL�z!V�RgW���m,M,c
U2|-E�����	�1U�$!U�sŗ�tr�KwK�+�6�Ϸ���ې�cdF'�G��O[$MwiOȫ̬ʴLC�ph���t{"W�""BAy?��^����E/샳%�B�6��=<�	N�=O-�CtJcȉI�+P�n{�{�V��^SI��.��֍3��m�U+"���,5�	N�98o;ɯ,������#��U]��k�h:�2�Vr���^�uO����*�T�R��ˏ_��M� ����\Dzo��E�U�p7jѢ�D�Y�B�g����^��D�J��fO�u����]{"�a�ܴB�~H���MH��jI��뤣آN��4Us�b�f��`��9?4������W��m��4ʇz"�2�����bi�
U5t�9>_��*�b�&h�W��nzR.�:�4D���?F�!�ԛ�V��yo��ĵ/1��$}B����<o�}|�m��:�
�t�Ħ�mJ���b*��O�|��Ut,n�#�?Y���	�L�ɯG&�9�YM~��6�cv�@�B�����z���� ��f�c{��m��Ͷ��170�j�}�OD��O��o\�MplmS�.�勬�o���P6��'{yox�{������(��Z�.�u�z�s?Qd��TW[�N�������p�Bp�q�W��Tv�H/�m�����D22�9ѵ����&Q�X�mBoFs�X��*J ��^I�23ۀ���P��8�z%&��@�\�o���]�_� x�&��G���i�����J6*�w!���1���ә>R�޼mbK��:m�]>�Ҍ^4��:_#	��tC.�����P�db%�*��5���ǥ�`%��B�7�����c�ۯ�̭_?Q�]ŗR� ]���xP����B�߫z"�ˬ"mL����~T�MwII\����9�n^���?F��� ��ݙ�o1�VN�V�6>�B��m��������&�3'5��k�i�왕���4)vmH�
3)���Z�5�g�F�2���+)�+�Ӊ|�3�o8e�Z-�3p���s6J�#&�z�ٖ�B>f�֏�u��gI>fI�SS� ��u&�(�N���s��M��|{�	��HW��_����a�<��0�>w)F)�g��B5�xw|�&�������M�rV:�~O�iv̜�N�;��I	�(E��bTp��p_=��z�iJ���]lؑ��޳�V7�k�����{��#��� '�mJ���F��`�`1؃ׇ7ח���R:��;v�Z�Ab4k�=��6�3�w�~"�L���/�y�f67���ÂB�+&9���{S9�B��{]+3bq��1B�xC�ߏ�cx�˺�ٺ���X
t�
�ܺ��uJJ��L���QyQ�mr.W�*\9��}2��(2�n�w��ݙ
��vcG�_7ڑʿ���D��̢X�U�+I�����_��S�|9�Nd�3J���
~����Z����� a*�$����[(�����$],�~:ř��~|rِ@��O�%Il%�����C�EJ&��B���NBx�)�VS]�DKi~��c(m~�� �Ĉ�9q+'b�$'��ن�-`�	�����d����yS�ǚ�S@�ʽ��c=}S,PB(�5&�^]��1v�_u&���dd�I�i���Ӻ·$!�d�.�q�.�j.���,ۨ�d�U��C�Q��?�q3�Zo`r�0��/�����|��)M��t\��B�c$�.Q.ͦ�d�6i�z|r��<��-څ�-j�~�fe�VUxs�S{B]c�����������\�G��#�1���3�����H#���7F+�=�Lʲ�jl��/�572��\�.7�N������!�ZD[[�?Jw%�'_�!��)0)���>Sb�䎒bJ�����)O&�I�
��c�WrG���,�i^Jh1C�I(�bQ7!�|�F��Z�*h��5��n�����}���w
6K�����s��i�@�'�߽�_�\����'�DQ��D�K�I�JD�xI�<�~4�F��=�7O֑��l{�B�PO;;vdD�,���5�%(v�HapL�M�8�Z��\�}������!����xy<M�R������a�������"*
	X�оNLN~B{��x%��Ww��7pt��(���8
��(`���	��y!7����{�O�~��ǋD��K���멽���$Sin���]��Ck͇�cJ�6� L���rA��c,т}Q�9;�����2�\��t�+���?1��e7/'�����fTr�1����tJ����iE���8�{f���v�]1���c�5��9�)��"\��GıL�'�m������]�M��d�w���{�nO�I�p���d>�������:r�f��1���քK�Nn�ԉ�)�UCib�����,�/��1�Bsw\뉬��%�$AX�V!���cʗa��| �Q�ѯ�!��/)���W|�����L��� ]��w�uO��yWz#�Ƚ����v��VF̊�N��� Z����G�y�X ����g�lX�&O�HR�:p:�ݻ@���O�R�e>rj��)��?���G������*��"��h7�>���R􊨷��/�~��d�UЯ��D��B�Vx�@�G�ٝ��
�@.��]���Lv�Dl��{,,�%������G�!�B�~+I�`���S�wg���uvٸ*������ڃ��9m�he�wL����O'�N��HT�A��8��죞�{�!t�������!k4n9?���,���Z3�À�_�}Ԝ��U��o�?�H�!��$���x��-m��A?�"�ݟ�+ʪɔJ���PK   ���X}�  �*     jsons/user_defined.json�Zio�H�+�>�b�D߇�)�쎱�m��.�0�>2�PR2F���Eɲc�P�60��'�ǫbw��zE~�,�n��`�Z��7bY?�N��fQ���9�	Y�������߷��؛����!;k�L��dg��Y�Ue3������Epv>�� L.�\vto�z:)=�of#�C<h��5
q�
/	q������P-��N����-���Y�����5��r�8�OrV:�?X�Y�т�%F2\Y$=���@���m�	�+]]��$9�(��X�5e���@ʺ���u4d{Ӎ������s�9��Y�9��۲:�b=9�>�V7G��vn��9���k�%\�x�c�m}��Xh�7�=YU�<Uu�ϗM	�a���E��P��5f4g�k>���D���Ŭr���ޮ�������p�c�Oz�Yα�r��ʥd�<��v��	����b� ��c,�TI�a���.>�9Sʨ)5&'L(��_'G��델�p�[�@��CM}�e�f�u��S���*�:�<9}Ə�kj��eS��i)�$��}Xӆ2_�RB w8v���`pD	�9�$�!r�51����WH� ��T8��#;~)Z�y���9XU����&}M����������<�<��h�&��ٶ�~��{.I��",��W"�`YήQyU%��aL���I�k:��.�y5��R�zǆ@u�&��� ��b0�9&�.�hZ���0h�T4-�gl�K)��3>�%M�����<�x'����a�F�Dأ�0l�H�l,�.�M�#+���4�#2\]n�
;L�S�D*�0iiOђ������-�k�Q{j�ND�è]���v
�F�r��DT9�ڥغ��g�S�X"�pB�=��'�Ӌ��.��:�.�S�d"�0�XO�R��xH<JG'��Q��7uD� E���3��'���V�/6�B��7�U���|�V�Gm���-�������T�ǭ��*e1ǚ�e��w�@��3d�V�h�rՀ0���F�����?��{ĕ��Y�����{F����f�lS�x$��5a����f���\�<��7��}��<T��y�̶���"9�Eo-r�Z�	H`�u��H�d�&�GH0�
n@��¦��X�aØ�R����/�*���=��;�~�cl�0"�{j�n�=:���qo����$׭slo�'���[��K��n�{ka�uP����;�����Qa�D<(�4����r,1�H�п�?$�n3�q�W�=���.۾?>gG�f����~/�̹0�^�N�Jy1��³1K<��XXn�J�F/#�4�Di�) J���C�MI��������t�i	��|�|*���0z�l���f7�D&�ώG�n���l��S�1��>�+B���7`��V�a�` 5������q�R�G'�]���oQ����1Hߢ����Y�WIK�=&�7)�=s5H�$g��/A��5L�ff�3x��(ΕQx�k���P=�,h0���g��o8���Я�&��Ȝs#4|�c��wi���3/��3�s,�صˣ{�39x�'��I��kv�g��ŧ��X�� k��'��K����/���AG��R2��%��BC/u�k9ϝ+7h��wESg��Y܆���w�7Qi�\dH����AZ� �*�8K�ç7�f�Bv�
�?�E��ГbΑ %����yX�����۶���wz2^��+�pB;�^�̀�%����T�|�kVL�Ph)�fT�hJG�\� ��q������b�	�)�>�%���dў���w���(�=y�<�=��f�;�)u�}�W��M��o;>���y� "#��)�$�XD�
ɌK�SR�ȵAL�8�0H��R��{���V�> 
��f��B��� S\�B��W��2v�h�m�g����w �$�rhPT�v�C�_gڠ��}r�;�(7�]!\�h��_�\8:�z�7�W�ֈ�VD��Q��K���q���j�O�F�7����C���o?L#�@�`K�9nm��0J�T�� q��!�@ׂ#�wB)w�H&b��C<��8�8y�g(pɘ��ߎ��6�{��`�I���n��a�(�_�u4Z{A�B!�Z�ȑ� 8
�!�S�������PK
   ���X_d�y  H�                   cirkitFile.jsonPK
   ���Xx�آ  �  /             �  images/0fa89018-bbd7-413a-af56-bcf37033748d.pngPK
   ���X��<�8� � /             �.  images/20128c01-dfdf-4258-b49d-382729dffbb1.pngPK
   9l�X�o��  �  /              images/54b474af-19f8-4da8-b85c-ecb600c58ca3.pngPK
   ���X�\�]�� �� /             �4 images/8e60f633-70d2-40b4-a331-b1224c91635f.pngPK
   ���X���<  -  /             � images/988d5287-ee6b-46f4-9561-988eb80bd729.pngPK
   9l�X�� �  �  /             d3 images/a80855a5-8bca-4bf2-b044-5bb17264cccb.pngPK
   ���X���8  8  /             IQ images/c52c1984-b936-4e70-81fd-2ef40f9d3319.pngPK
   ���X$7h�!  �!  /             �� images/c6364832-c854-438f-b38b-75bf2a0cd33f.pngPK
   ���XGJ���0  �0  /             � images/cfd0a77b-9a45-4601-b836-f8aa27cd4ccb.pngPK
   ���X��k�  n /             �� images/e6413bd2-a01a-4823-b22b-7acb31e08f91.pngPK
   ���XKm���[ � /             (� images/e677f489-379d-40e3-bb59-6fe87b8e7dd0.pngPK
   ���X��6�  S# /             @: images/ea543ea3-2b47-4327-947a-6d32920e175d.pngPK
   ���XF1��^$ �B /             �[ images/efd6e310-ffe8-4178-823b-653710540121.pngPK
   ���XP��/�  ǽ  /             5� images/f42d805d-3c79-4d19-85d7-77e6ec425ca7.pngPK
   ���X}�  �*               �2 jsons/user_defined.jsonPK      �  F;   